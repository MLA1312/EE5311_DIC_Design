** sch_path: /home/EE23B038/ee5311/tutorial_2/tutorial_2_1a.sch
**.subckt tutorial_2_1a
XM1 Vin Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vin Vin GND 1.8
**** begin user architecture code

.control
dc Vin 0 1.8 0.01
let mu = 0.025
let WbyL = 0.42/0.15
let Cox = 0.00834
let Vth = 0.7
let vsat = 8e4
let Vgs = V(Vin)
let Vds = Vgs
let lamban = 0.2
let Ecl = 2*vsat * 0.15e-6/mu
let Vgt = max(Vgs-Vth,0)
let Vdsat = (Vgt)*Ecl/(Vgt + Ecl)
let Vmin = min(Vgs, Vdsat)
let idfit = 0.5*mu*Cox*WbyL*Ecl*(Vgt^2)*(1+lamban*Vds)/(Vgt+Ecl)
set filetype=ascii
wrdata nmos_ids_vgs.txt -I(Vin) idfit
plot -I(Vin) idfit
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
