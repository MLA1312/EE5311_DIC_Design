** sch_path: /home/global/EE23B038/tutorial_6/6.1v2/inv.sch
.subckt inv DVDD in out DGND
*.PININFO in:I DVDD:B DGND:B out:O
XM1 out in DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 out in DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM3 net1 out DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 net1 out DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
.ends
.end
