** sch_path: /home/EE23B038/ee5311/tutorial_2/tutorial_2_1b.sch
**.subckt tutorial_2_1b
XM1 net1 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdd1 net1 GND 1.8
Vin1 net2 GND 1.8
**** begin user architecture code

.control
let Vgs = 0.6
let mu = 0.025
let WbyL = 0.42/0.15
let Cox = 0.00834
let Vth = 0.7
let vsat = 8e4
let lambdan = 0.2
let EcL = 2*vsat* 0.15e-6/mu
repeat 4
  alter Vin1 $&Vgs
  dc Vdd1 0 1.8 0.02
  let Vds = "v-sweep"
  let Vds1 = min(Vgs - Vth, Vds)
  let Vgt = max(Vgs - Vth, 0)
  let Vds_min = min(Vds1, EcL*Vgt/(EcL+Vgt))
  let idfit = mu*Cox*WbyL*EcL*(Vgs - Vth - Vds_min / 2)*Vds_min*(1 + lambdan * Vds)/(Vgt + EcL)
  let Vgs = Vgs + 0.4
end
plot dc1.I(Vdd1)*-1 dc2.I(Vdd1)*-1 dc3.I(Vdd1)*-1 dc4.I(Vdd1)*-1 dc1.idfit dc2.idfit dc3.idfit dc4.idfit
set filetype=ascii
wrdata nmos_ids_vds.txt dc1.I(Vdd1)*-1 dc2.I(Vdd1)*-1 dc3.I(Vdd1)*-1 dc4.I(Vdd1)*-1 dc1.idfit dc2.idfit dc3.idfit dc4.idfit
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
