** sch_path: /home/EE23B038/ee5311/tutorial_3/tutorial_3_1a.sch
**.subckt tutorial_3_1a
XM1 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vin1 Vin GND 1.8
Vdd1 VDD GND 1.8
**** begin user architecture code


.control
dc Vin1 0 1.8 0.01
plot v(Vout) v(Vin)
let derivout = deriv(v(Vout))
plot derivout
meas dc Vil when derivout=-1 cross=1
meas dc Vih when derivout=-1 cross=2
meas dc Vm when v(Vout)=0.9
let NMl=Vil
let NMh=1.8 - Vih
echo NML: $&NMl NML: $&NMh
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
