** sch_path: /home/global/EE23B038/tutorial_7/tutorial_7v2.sch
**.subckt tutorial_7v2
Vin1 Vin GND PULSE(0 1.8 10ps 5ps 5ps 200ps 400ps)
Vdd1 VDD GND 1.8
x1 VDD Vout Vin GND nors
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.include nors_extracted.spice
.control
tran 0.01p 400p
plot v(Vout) v(Vin)
meas tran thl trig v(Vin) val=0.9 rise=1 targ v(Vout) val=0.9 fall=1
meas tran tlh trig v(Vin) val=0.9 fall=1 targ v(Vout) val=0.9 rise=1
let delay = ( $&thl + $&tlh ) / 2
echo delay : $&delay
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
