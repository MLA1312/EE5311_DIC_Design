* NGSPICE file created from fa16.ext - technology: sky130A

.subckt fa16 S15 DVDD A12 A13 A14 A15 A9 A8 A10 A11 B13 B12 A6 B14 A5 A4 B15 A7 A2 B11 B10 A0 B9 B8 A1 A3 B6 B5 B4 B7 B2 B0 B3 B1
+ Cin DGND
X0 a_4691_n3974# A11.t0 DGND.t285 DGND.t284 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_5402_n3546# a_4204_n3054# a_5819_n3308# DVDD.t272 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_4691_n1494# A15.t0 DGND.t390 DGND.t389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_541_n828# A2.t0 DVDD.t107 DVDD.t106 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 DVDD.t507 a_1201_n3054# a_2273_n2734# DVDD.t506 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X5 a_5288_n828# B14.t0 a_5192_n828# DVDD.t232 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 DGND.t541 B9.t0 a_4363_n2434# DGND.t540 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_4697_n2434# B9.t1 a_3946_n2306# DGND.t344 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_894_n1194# a_143_n1036# a_798_n1194# DGND.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 DGND.t160 A10.t0 a_5456_n3674# DGND.t159 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X10 a_894_n3674# a_143_n3516# a_798_n3674# DGND.t211 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 DGND.t340 A14.t0 a_5456_n1194# DGND.t339 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X12 DVDD.t109 A2.t1 a_n41_n1814# DVDD.t108 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_n131_n574# a_n71_n600# DGND.t528 DGND.t527 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X14 a_1467_46# A1.t0 DGND.t415 DGND.t414 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X15 a_4691_n1814# A15.t1 DVDD.t341 DVDD.t340 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 DVDD.t103 A6.t0 a_185_n3308# DVDD.t102 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_11_n1194# A2.t2 DGND.t468 DGND.t467 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X18 a_3874_n3700# a_5402_n3546# DGND.t238 DGND.t237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_11_n3674# A6.t1 DGND.t36 DGND.t35 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X20 a_3874_n1220# a_5402_n1066# DGND.t526 DGND.t525 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_5819_n2068# A8.t0 DVDD.t169 DVDD.t168 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 DVDD.t199 a_3861_n3080# a_3322_n4062# DVDD.t198 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X23 a_147_n1494# B2.t0 a_n131_n1814# DGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X24 a_147_n3974# B6.t0 a_n131_n4294# DGND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X25 a_315_n3054# A4.t0 DVDD.t116 DVDD.t115 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 DGND.t10 B2.t1 a_n71_n1840# DGND.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 DGND.t183 B6.t1 a_n71_n4320# DGND.t182 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_3832_46# B13.t0 a_3736_46# DGND.t473 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_3655_n1516# a_3322_n1582# DVDD.t449 DVDD.t448 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_966_n3674# B6.t2 a_894_n3674# DGND.t472 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 a_4523_n3054# B9.t2 a_4441_n3054# DVDD.t514 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_2350_46# a_636_n574# a_2254_46# DGND.t151 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_3874_20# a_5402_174# DGND.t351 DGND.t350 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X34 a_966_n1194# B2.t2 a_894_n1194# DGND.t416 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X35 DGND.t283 A11.t1 a_4441_n4294# DGND.t282 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 DGND.t343 A15.t2 a_4441_n1814# DGND.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 a_3765_n3080# a_4441_n3054# a_4691_n3054# DVDD.t490 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X38 DVDD.t15 B10.t0 a_5456_n3308# DVDD.t14 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 a_3736_n3308# A11.t2 DVDD.t286 DVDD.t285 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X40 a_3874_n1220# a_5402_n1066# DVDD.t530 DVDD.t529 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X41 DVDD.t154 A13.t0 a_4523_n574# DVDD.t153 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X42 a_5192_n1194# A14.t1 DGND.t496 DGND.t495 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X43 a_5192_n3674# A10.t1 DGND.t273 DGND.t272 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X44 DVDD.t216 a_1557_n2434# a_143_n3516# DVDD.t215 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X45 a_2273_n254# a_1201_n1814# DVDD.t305 DVDD.t304 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 a_n71_n600# B0.t0 a_315_n574# DVDD.t6 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X47 DGND.t185 A7.t0 a_1641_n3674# DGND.t184 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X48 a_6153_n2068# B8.t0 a_5402_n2306# DVDD.t312 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X49 a_n41_n1814# B2.t3 DVDD.t409 DVDD.t408 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X50 DGND.t440 A3.t0 a_1641_n1194# DGND.t439 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X51 a_n41_n1814# a_n71_n1840# a_n131_n1814# DVDD.t42 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X52 a_1641_412# a_636_n574# a_1557_46# DVDD.t145 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X53 a_5819_n828# A14.t2 DVDD.t495 DVDD.t494 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X54 a_n71_n1840# B2.t4 a_315_n1814# DVDD.t381 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X55 a_3765_n3080# B9.t3 a_4691_n2734# DGND.t512 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X56 DVDD.t227 A15.t3 a_4523_n1814# DVDD.t226 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X57 a_4697_n828# B15.t0 a_3946_n1066# DVDD.t247 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X58 a_11_46# A0.t0 DGND.t72 DGND.t71 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X59 a_5360_n2434# a_2995_n4294# a_5288_n2434# DGND.t61 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X60 a_541_n828# B2.t5 DVDD.t364 DVDD.t363 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X61 DVDD.t274 A10.t2 a_5855_n4294# DVDD.t273 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X62 DVDD.t537 A0.t1 a_185_412# DVDD.t536 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X63 DVDD.t175 A13.t1 a_4697_412# DVDD.t174 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X64 a_1641_n2434# a_636_n3054# a_1557_n2434# DGND.t142 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 a_4000_n2068# a_3946_n2306# a_3904_n2434# DVDD.t323 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 DVDD.t293 B12.t0 a_6023_n574# DVDD.t292 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X67 a_894_n828# a_143_n1036# a_798_n1194# DVDD.t3 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_2422_n2434# B5.t0 a_2350_n2434# DGND.t307 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X69 a_185_n2068# B4.t0 DVDD.t183 DVDD.t182 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X70 a_3655_n3996# a_3322_n4062# DVDD.t193 DVDD.t192 sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 DVDD.t139 A10.t3 a_6153_n3308# DVDD.t138 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X72 DVDD.t303 a_2908_n600# S15.t1 DVDD.t302 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X73 a_3655_n3996# a_3322_n4062# DGND.t199 DGND.t198 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X74 a_3655_n1516# a_3322_n1582# DGND.t457 DGND.t456 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X75 a_4000_46# a_3946_174# a_3904_46# DGND.t356 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_1467_n1194# A3.t1 DGND.t113 DGND.t112 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X77 a_1467_n3674# A7.t1 DGND.t386 DGND.t385 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X78 a_5456_n3308# a_4204_n3054# DVDD.t271 DVDD.t270 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X79 DVDD.t311 A12.t0 a_5456_412# DVDD.t310 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X80 a_1201_n3054# a_1261_n3080# DGND.t221 DGND.t220 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X81 DVDD.t133 a_636_n3054# a_1997_n2068# DVDD.t132 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X82 a_5402_n2306# a_2995_n4294# a_5819_n2068# DVDD.t50 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X83 a_101_n2434# B4.t1 a_11_n2068# DVDD.t423 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X84 DGND.t464 B11.t0 a_4363_n3674# DGND.t463 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 DGND.t494 A0.t2 a_185_46# DGND.t493 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X86 a_4363_46# A13.t2 DGND.t40 DGND.t39 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X87 DGND.t120 B15.t1 a_4363_n1194# DGND.t119 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X88 a_4697_n1194# B15.t2 a_3946_n1066# DGND.t97 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X89 a_4697_n3674# B11.t1 a_3946_n3546# DGND.t465 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 a_4697_412# B13.t1 a_3946_174# DVDD.t75 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X91 DGND.t219 a_143_n2276# a_541_n2434# DGND.t218 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X92 DVDD.t229 A15.t4 a_4697_n828# DVDD.t228 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X93 a_1557_n2434# B5.t1 a_1467_n2434# DGND.t186 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X94 DVDD.t250 a_3669_n342# a_3322_n1582# DVDD.t249 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 a_2790_n3928# a_1968_n4294# a_2569_n4255# DGND.t466 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X96 a_798_n3674# a_101_n3674# a_541_n3308# DVDD.t26 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X97 a_1641_n2434# B5.t2 DGND.t297 DGND.t296 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X98 a_2790_n1448# a_1968_n1814# a_2569_n1775# DGND.t54 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X99 DVDD.t288 A0.t3 a_n41_n574# DVDD.t287 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X100 a_4000_n2434# a_3874_n2460# DGND.t260 DGND.t259 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 DVDD.t466 A4.t1 a_185_n2068# DVDD.t465 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X102 a_3543_n342# a_5773_n1814# a_6023_n1814# DVDD.t170 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X103 a_4697_46# B13.t2 a_3946_174# DGND.t480 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X104 a_6023_n254# A12.t1 DGND.t13 DGND.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 a_2908_n600# a_3874_n1220# a_3832_n828# DVDD.t127 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X106 a_4363_n828# A15.t5 DVDD.t475 DVDD.t474 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X107 a_3736_46# A13.t3 DGND.t85 DGND.t84 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X108 a_185_412# Cin.t0 a_101_46# DVDD.t496 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X109 a_3832_n3308# B11.t2 a_3736_n3308# DVDD.t37 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X110 a_1997_n3308# B7.t0 DVDD.t414 DVDD.t413 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X111 DGND.t99 A9.t0 a_4697_n2434# DGND.t98 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X112 a_315_n4294# A6.t2 DVDD.t122 DVDD.t121 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X113 a_2254_46# a_1557_46# a_1997_46# DGND.t235 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X114 DGND.t373 A5.t0 a_1479_n2734# DGND.t372 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X115 a_101_n1194# B2.t6 a_11_n828# DVDD.t435 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X116 DVDD.t459 A2.t3 a_185_n828# DVDD.t458 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X117 a_3946_n3546# a_3874_n3700# a_4363_n3308# DVDD.t487 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 a_4523_n4294# B11.t3 a_4441_n4294# DVDD.t7 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X119 DGND.t174 a_5773_n574# a_3861_n600# DGND.t173 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X120 a_3669_n2822# a_4441_n4294# a_4691_n4294# DVDD.t358 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X121 DVDD.t462 a_1557_n3674# a_1968_n4294# DVDD.t461 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X122 DVDD.t236 B8.t1 a_5456_n2068# DVDD.t235 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 a_3736_n2068# A9.t1 DVDD.t360 DVDD.t359 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X124 a_1557_46# B1.t0 a_1467_412# DVDD.t535 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X125 DVDD.t189 A4.t2 a_n41_n3054# DVDD.t188 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X126 DGND.t488 a_4441_n3054# a_3765_n3080# DGND.t487 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X127 a_4204_n3054# a_3946_n2306# DGND.t324 DGND.t323 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X128 a_1997_n3308# A7.t2 DVDD.t443 DVDD.t442 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X129 a_4691_n3054# A9.t2 DVDD.t173 DVDD.t172 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X130 a_3669_n2822# B11.t4 a_4691_n3974# DGND.t462 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X131 DGND.t407 a_5773_n3054# a_3861_n3080# DGND.t406 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X132 a_3669_n342# B15.t3 a_4691_n1494# DGND.t25 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X133 a_2459_n254# a_1201_n574# a_2363_n254# DGND.t143 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X134 a_2254_n1194# a_1557_n1194# a_1997_n828# DVDD.t398 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X135 DGND.t516 A9.t3 a_4000_n2434# DGND.t515 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X136 a_3946_174# a_3874_20# a_4363_412# DVDD.t268 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_5360_n1194# a_4204_n574# a_5288_n1194# DGND.t207 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X138 a_5360_n3674# a_4204_n3054# a_5288_n3674# DGND.t271 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X139 a_1641_n3674# a_636_n4294# a_1557_n3674# DGND.t31 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 DVDD.t464 A6.t3 a_966_n3308# DVDD.t463 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X141 DGND.t109 B1.t1 a_1261_n600# DGND.t108 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 a_3795_n254# a_3765_n600# a_3711_n254# DGND.t400 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X143 a_1641_n1194# a_636_n1814# a_1557_n1194# DGND.t252 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X144 a_2422_n1194# B3.t0 a_2350_n1194# DGND.t241 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X145 a_2422_n3674# B7.t1 a_2350_n3674# DGND.t335 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X146 a_4000_46# a_3874_20# DGND.t267 DGND.t266 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X147 DVDD.t30 A8.t1 a_6153_n2068# DVDD.t29 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X148 a_1479_n2734# B5.t3 a_1201_n3054# DGND.t306 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X149 a_4363_n3308# A11.t3 DVDD.t284 DVDD.t283 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X150 a_3904_46# a_3874_20# a_3832_46# DGND.t265 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X151 DVDD.t77 B15.t4 a_4691_n1814# DVDD.t76 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X152 a_1467_412# A1.t1 DVDD.t429 DVDD.t428 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X153 DGND.t287 A0.t4 a_966_46# DGND.t286 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X154 a_3874_n2460# a_5402_n2306# DVDD.t196 DVDD.t195 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X155 a_2422_46# B1.t2 a_2350_46# DGND.t163 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X156 a_5456_n2068# a_2995_n4294# DVDD.t49 DVDD.t48 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X157 a_1201_n1814# a_1261_n1840# DGND.t428 DGND.t427 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X158 a_1201_n4294# a_1261_n4320# DGND.t380 DGND.t379 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X159 a_966_n828# B2.t7 a_894_n828# DVDD.t12 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 a_n41_n3054# B4.t2 DVDD.t387 DVDD.t386 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X161 a_n41_n3054# a_n71_n3080# a_n131_n3054# DVDD.t313 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X162 a_11_n828# A2.t4 DVDD.t318 DVDD.t317 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X163 DVDD.t493 A14.t3 a_5456_n828# DVDD.t492 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X164 a_n71_n3080# B4.t3 a_315_n3054# DVDD.t159 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X165 a_5855_n574# B12.t1 a_5773_n574# DVDD.t18 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X166 DVDD.t164 B15.t5 a_4000_n828# DVDD.t163 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 DVDD.t141 A10.t4 a_5456_n3308# DVDD.t140 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X168 a_894_n3308# a_143_n3516# a_798_n3674# DVDD.t213 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X169 DVDD.t343 A9.t4 a_4523_n3054# DVDD.t342 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 DVDD.t451 a_3861_n600# a_3322_n1582# DVDD.t450 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X171 DGND.t210 a_143_n3516# a_541_n3674# DGND.t209 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X172 DGND.t2 a_143_n1036# a_541_n1194# DGND.t1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 a_6023_n2734# A8.t2 DGND.t79 DGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X174 a_6153_46# B12.t2 a_5402_174# DGND.t290 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X175 a_1557_n3674# B7.t2 a_1467_n3674# DGND.t367 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X176 a_1557_n1194# B3.t1 a_1467_n1194# DGND.t384 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X177 a_798_n2434# a_101_n2434# a_541_n2068# DVDD.t316 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X178 a_1641_n1194# B3.t2 DGND.t509 DGND.t508 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X179 a_1641_n3674# B7.t3 DGND.t294 DGND.t293 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 a_2497_n1775# a_2315_n1775# DVDD.t353 DVDD.t352 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X181 a_4000_n1194# a_3874_n1220# DGND.t135 DGND.t134 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X182 a_4000_n3674# a_3874_n3700# DGND.t484 DGND.t483 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X183 a_11_n3308# A6.t4 DVDD.t64 DVDD.t63 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X184 a_541_412# B0.t1 DVDD.t71 DVDD.t70 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 a_541_n2434# B4.t4 DGND.t311 DGND.t310 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X186 a_1997_46# B1.t3 DGND.t292 DGND.t291 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X187 DVDD.t327 a_3226_n4062# a_3177_n4294.t1 DVDD.t326 sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X188 DGND.t477 A15.t6 a_4697_n1194# DGND.t476 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X189 DGND.t281 A11.t4 a_4697_n3674# DGND.t280 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X190 a_3832_n2068# B9.t4 a_3736_n2068# DVDD.t328 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X191 a_1997_n2068# B5.t4 DVDD.t181 DVDD.t180 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X192 DGND.t426 A1.t2 a_1479_n254# DGND.t425 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X193 a_3627_n254# a_3543_n342# DGND.t137 DGND.t136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X194 a_541_46# B0.t2 DGND.t168 DGND.t167 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X195 DGND.t27 A12.t2 a_5456_46# DGND.t26 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X196 a_147_n254# B0.t3 a_n131_n574# DGND.t166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X197 DGND.t438 A3.t2 a_1479_n1494# DGND.t437 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X198 DGND.t388 A7.t3 a_1479_n3974# DGND.t387 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X199 a_966_n3308# B6.t3 a_894_n3308# DVDD.t483 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X200 a_2254_n2434# a_1557_n2434# a_1997_n2434# DGND.t214 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X201 a_2350_412# a_636_n574# a_2254_46# DVDD.t144 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X202 a_3946_n2306# a_3874_n2460# a_4363_n2068# DVDD.t261 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 a_5288_n2434# B8.t2 a_5192_n2434# DGND.t539 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X204 a_5192_n3308# A10.t5 DVDD.t99 DVDD.t98 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X205 a_1641_n828# B3.t3 DVDD.t325 DVDD.t324 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X206 a_2254_46# a_1557_46# a_1997_412# DVDD.t240 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X207 a_5360_46# a_3177_n4294.t2 a_5288_412# DVDD.t150 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X208 a_894_46# Cin.t1 a_798_46# DGND.t403 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X209 DVDD.t101 A6.t5 a_n41_n4294# DVDD.t100 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X210 DGND.t366 a_4441_n4294# a_3669_n2822# DGND.t365 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X211 DVDD.t441 A7.t4 a_1641_n3308# DVDD.t440 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X212 a_2569_n1775# a_1968_n1814# a_2497_n1775# DVDD.t43 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X213 a_3765_n600# a_4441_n574# a_4691_n574# DVDD.t137 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X214 DGND.t145 a_4441_n1814# a_3669_n342# DGND.t144 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X215 a_5192_46# A12.t3 DGND.t170 DGND.t169 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X216 DGND.t300 A12.t4 a_5773_n574# DGND.t299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X217 a_798_n1194# a_101_n1194# a_541_n828# DVDD.t375 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X218 a_2497_n4255# a_2315_n4255# DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_3434_n4026# a_3946_n3546# DGND.t263 DGND.t262 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X220 DGND.t418 B5.t5 a_1261_n3080# DGND.t417 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X221 a_1997_n2068# A5.t1 DVDD.t334 DVDD.t333 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X222 a_3434_n1546# a_3946_n1066# DGND.t116 DGND.t115 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X223 a_4691_n4294# A11.t5 DVDD.t282 DVDD.t281 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X224 DVDD.t105 A3.t3 a_1291_n1814# DVDD.t104 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X225 a_3874_20# a_5402_174# DVDD.t348 DVDD.t347 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X226 DGND.t256 a_5773_n4294# a_3543_n2822# DGND.t255 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X227 a_3861_n3080# a_5773_n3054# a_6023_n3054# DVDD.t407 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X228 DGND.t172 a_5773_n1814# a_3543_n342# DGND.t171 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X229 a_4363_412# A13.t4 DVDD.t36 DVDD.t35 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X230 DGND.t150 a_636_n574# a_1997_46# DGND.t149 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X231 DGND.t254 A15.t7 a_4000_n1194# DGND.t253 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X232 DGND.t279 A11.t6 a_4000_n3674# DGND.t278 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X233 DVDD.t437 A4.t3 a_966_n2068# DVDD.t436 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X234 DVDD.t256 A15.t8 a_4000_n828# DVDD.t255 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X235 a_2363_n2734# a_n131_n3054# a_2273_n2734# DGND.t474 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X236 a_5456_412# a_5402_174# a_5360_46# DVDD.t346 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X237 a_5360_46# a_3177_n4294.t3 a_5288_46# DGND.t511 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X238 a_6153_n828# B14.t1 a_5402_n1066# DVDD.t532 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X239 a_541_n2434# A4.t4 DGND.t536 DGND.t535 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X240 a_1479_n1494# B3.t4 a_1201_n1814# DGND.t73 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X241 a_1479_n3974# B7.t4 a_1201_n4294# DGND.t175 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X242 a_3434_n1546# a_3946_n1066# DVDD.t112 DVDD.t111 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X243 a_3861_n3080# B8.t3 a_6023_n2734# DGND.t96 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X244 a_4363_n2068# A9.t5 DVDD.t57 DVDD.t56 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X245 a_1467_n3308# A7.t5 DVDD.t389 DVDD.t388 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X246 DGND.t328 B9.t5 a_4000_n2434# DGND.t327 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 a_3874_n3700# a_5402_n3546# DVDD.t243 DVDD.t242 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X248 DVDD.t209 B13.t3 a_4000_412# DVDD.t208 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 DGND.t243 B12.t3 a_5456_46# DGND.t242 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X250 a_2569_n4255# a_1968_n4294# a_2497_n4255# DVDD.t457 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X251 a_n41_n4294# a_n71_n4320# a_n131_n4294# DVDD.t491 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X252 a_n41_n4294# B6.t4 DVDD.t482 DVDD.t481 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X253 DGND.t22 B8.t4 a_5819_n2434# DGND.t21 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X254 a_n71_n4320# B6.t5 a_315_n4294# DVDD.t519 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X255 a_2569_n1448# a_2315_n1775# DGND.t358 DGND.t357 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X256 a_2569_n3928# a_2315_n4255# DGND.t5 DGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X257 DVDD.t454 B11.t5 a_4363_n3308# DVDD.t453 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X258 a_4697_n3308# B11.t6 a_3946_n3546# DVDD.t452 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X259 a_1261_n3080# A5.t2 DGND.t338 DGND.t337 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 DVDD.t280 A11.t7 a_4523_n4294# DVDD.t279 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X261 a_n131_n3054# a_n71_n3080# DGND.t315 DGND.t314 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X262 a_894_n2068# a_143_n2276# a_798_n2434# DVDD.t221 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X263 a_1291_n1814# B3.t5 DVDD.t205 DVDD.t204 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X264 a_1641_46# a_636_n574# a_1557_46# DGND.t148 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X265 DVDD.t11 A8.t3 a_5456_n2068# DVDD.t10 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X266 a_2422_n828# B3.t6 a_2350_n828# DVDD.t187 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X267 DGND.t453 a_n131_n1814# a_2543_n254# DGND.t452 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X268 a_6023_n3974# A10.t6 DGND.t107 DGND.t106 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X269 a_6023_n1494# A14.t4 DGND.t492 DGND.t491 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X270 a_4691_n254# A13.t5 DGND.t436 DGND.t435 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 a_1641_n828# a_636_n1814# a_1557_n1194# DVDD.t254 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X272 a_11_n2068# A4.t5 DVDD.t521 DVDD.t520 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X273 DVDD.t471 A14.t5 a_6153_n828# DVDD.t470 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X274 DVDD.t523 B9.t6 a_4691_n3054# DVDD.t522 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X275 a_2350_n2434# a_636_n3054# a_2254_n2434# DGND.t141 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X276 a_541_n1194# B2.t8 DGND.t442 DGND.t441 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X277 a_541_n3674# B6.t6 DGND.t118 DGND.t117 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X278 a_6023_n1814# A14.t6 DVDD.t473 DVDD.t472 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X279 DVDD.t309 A12.t5 a_6153_412# DVDD.t308 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X280 a_5360_n1194# a_4204_n574# a_5288_n828# DVDD.t203 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X281 a_2254_n1194# a_1557_n1194# a_1997_n1194# DGND.t399 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X282 a_2254_n3674# a_1557_n3674# a_1997_n3674# DGND.t471 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X283 a_966_n2068# B4.t5 a_894_n2068# DVDD.t406 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X284 DVDD.t534 B14.t2 a_5456_n828# DVDD.t533 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X285 a_5288_n1194# B14.t3 a_5192_n1194# DGND.t529 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X286 a_5288_n3674# B10.t1 a_5192_n3674# DGND.t100 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X287 a_3711_n2734# a_3669_n2822# a_3627_n2734# DGND.t222 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 a_5192_n2068# A8.t4 DVDD.t66 DVDD.t65 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X289 a_798_46# a_101_46# a_541_46# DGND.t95 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X290 a_3861_n600# a_5773_n574# a_6023_n574# DVDD.t171 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X291 a_3832_412# B13.t4 a_3736_412# DVDD.t467 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X292 a_6023_n574# A12.t6 DVDD.t395 DVDD.t394 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X293 a_4000_412# a_3874_20# DVDD.t267 DVDD.t266 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X294 DVDD.t114 A5.t3 a_1641_n2068# DVDD.t113 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X295 a_3736_412# A13.t6 DVDD.t34 DVDD.t33 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X296 a_2783_n1775# Cin.t2 a_2569_n1775# DVDD.t390 sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X297 DGND.t514 B7.t5 a_1261_n4320# DGND.t513 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X298 DGND.t7 B3.t7 a_1261_n1840# DGND.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X299 DGND.t434 A13.t7 a_4000_46# DGND.t433 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X300 a_3543_n2822# a_5773_n4294# a_6023_n4294# DVDD.t257 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X301 a_966_46# B0.t4 a_894_46# DGND.t138 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X302 a_5360_n3674# a_4204_n3054# a_5288_n3308# DVDD.t269 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X303 a_5456_n2434# a_5402_n2306# a_5360_n2434# DGND.t202 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X304 DVDD.t357 a_2273_n254# a_2783_n1775# DVDD.t356 sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X305 a_1641_n3308# a_636_n4294# a_1557_n3674# DVDD.t23 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X306 a_6153_412# B12.t4 a_5402_174# DVDD.t248 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 a_5773_n3054# B8.t5 DGND.t91 DGND.t90 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X308 DGND.t532 A5.t4 a_2422_n2434# DGND.t531 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X309 a_2422_n3308# B7.t6 a_2350_n3308# DVDD.t197 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X310 a_541_n1194# A2.t5 DGND.t320 DGND.t319 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X311 a_541_n3674# A6.t6 DGND.t195 DGND.t194 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X312 a_1291_n1814# a_1261_n1840# a_1201_n1814# DVDD.t434 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X313 a_966_412# B0.t5 a_894_412# DVDD.t405 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X314 DGND.t192 B13.t5 a_4000_46# DGND.t191 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_4441_n574# B13.t6 DGND.t538 DGND.t537 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_1261_n1840# B3.t8 a_1647_n1814# DVDD.t476 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X317 a_3543_n2822# B10.t2 a_6023_n3974# DGND.t105 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X318 a_3543_n342# B14.t4 a_6023_n1494# DGND.t530 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X319 a_n71_n600# A0.t5 DGND.t449 DGND.t448 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 DGND.t318 a_101_n2434# a_636_n3054# DGND.t317 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X321 DGND.t334 B15.t6 a_4000_n1194# DGND.t333 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X322 DGND.t460 B11.t7 a_4000_n3674# DGND.t459 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X323 a_1467_n2068# A5.t5 DVDD.t207 DVDD.t206 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X324 DVDD.t135 a_1201_n574# a_2273_n254# DVDD.t134 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X325 a_2569_n1775# Cin.t3 a_2569_n1448# DGND.t341 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X326 a_2569_n4255# a_143_n2276# a_2569_n3928# DGND.t217 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X327 a_3627_n2734# a_3543_n2822# DGND.t505 DGND.t504 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X328 a_185_n2434# a_143_n2276# a_101_n2434# DGND.t216 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_3322_n1582# a_3765_n600# DVDD.t400 DVDD.t399 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X330 DGND.t234 a_1557_46# a_143_n1036# DGND.t233 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X331 a_1261_n600# B1.t4 a_1647_n574# DVDD.t225 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X332 DGND.t486 B14.t5 a_5819_n1194# DGND.t485 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X333 DGND.t81 B10.t3 a_5819_n3674# DGND.t80 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X334 a_5402_174# a_3177_n4294.t4 a_5819_46# DGND.t70 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_2783_n4255# a_143_n2276# a_2569_n4255# DVDD.t220 sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X336 DVDD.t525 B9.t7 a_4363_n2068# DVDD.t524 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X337 a_5192_n828# A14.t7 DVDD.t345 DVDD.t344 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X338 a_1261_n4320# A7.t6 DGND.t44 DGND.t43 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X339 DVDD.t32 A5.t6 a_1291_n3054# DVDD.t31 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 a_n131_n1814# a_n71_n1840# DGND.t53 DGND.t52 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X341 a_1261_n1840# A3.t4 DGND.t503 DGND.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X342 a_n131_n4294# a_n71_n4320# DGND.t490 DGND.t489 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X343 a_4697_n2068# B9.t8 a_3946_n2306# DVDD.t290 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X344 DVDD.t489 B14.t6 a_6023_n1814# DVDD.t488 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X345 a_5192_412# A12.t7 DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X346 DGND.t302 a_n131_n4294# a_2543_n2734# DGND.t301 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X347 DVDD.t149 a_2273_n2734# a_2783_n4255# DVDD.t148 sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X348 DVDD.t212 a_143_n3516# a_541_n3308# DVDD.t211 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X349 a_1557_n3674# B7.t7 a_1467_n3308# DVDD.t401 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X350 DGND.t155 a_2273_n2734# a_2790_n3928# DGND.t154 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X351 DGND.t364 a_2273_n254# a_2790_n1448# DGND.t363 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X352 a_1641_n3308# B7.t8 DVDD.t339 DVDD.t338 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X353 a_4000_n3308# a_3874_n3700# DVDD.t486 DVDD.t485 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 a_3904_n2434# a_3874_n2460# a_3832_n2434# DGND.t258 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X355 a_4204_n3054# a_3946_n2306# DVDD.t322 DVDD.t321 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X356 a_2350_n3674# a_636_n4294# a_2254_n3674# DGND.t30 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X357 a_1647_n1814# A3.t5 DVDD.t86 DVDD.t85 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X358 a_2350_n1194# a_636_n1814# a_2254_n1194# DGND.t251 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X359 DVDD.t299 B11.t8 a_4691_n4294# DVDD.t298 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X360 a_5288_412# B12.t5 a_5192_412# DVDD.t123 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X361 DVDD.t278 A11.t8 a_4697_n3308# DVDD.t277 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X362 a_n41_n574# a_n71_n600# a_n131_n574# DVDD.t531 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X363 a_3226_n1582# a_3177_n4294.t5 a_3368_n1775# DVDD.t479 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X364 a_1997_412# A1.t3 DVDD.t427 DVDD.t426 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X365 DVDD.t433 A0.t6 a_966_412# DVDD.t432 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X366 a_4204_n574# a_3946_174# DGND.t355 DGND.t354 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X367 DVDD.t505 A13.t8 a_4000_412# DVDD.t504 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X368 a_1291_n3054# B5.t6 DVDD.t385 DVDD.t384 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X369 DVDD.t425 A1.t4 a_1291_n574# DVDD.t424 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X370 a_3322_n1582# a_3543_n342# DVDD.t129 DVDD.t128 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X371 a_n41_n574# B0.t6 DVDD.t368 DVDD.t367 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X372 DVDD.t253 a_636_n1814# a_1997_n828# DVDD.t252 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X373 a_5819_n2434# A8.t5 DGND.t111 DGND.t110 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X374 DVDD.t276 A11.t9 a_4000_n3308# DVDD.t275 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X375 a_5456_n1194# a_5402_n1066# a_5360_n1194# DGND.t524 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X376 a_5456_n3674# a_5402_n3546# a_5360_n3674# DGND.t236 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X377 a_5360_n2434# a_2995_n4294# a_5288_n2068# DVDD.t47 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X378 a_1997_46# A1.t5 DGND.t445 DGND.t444 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X379 a_5402_174# a_3177_n4294.t6 a_5819_412# DVDD.t410 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X380 a_1641_n2068# a_636_n3054# a_1557_n2434# DVDD.t131 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X381 a_5773_n4294# B10.t4 DGND.t232 DGND.t231 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X382 a_5773_n1814# B14.t7 DGND.t65 DGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X383 DGND.t346 Cin.t4 a_541_46# DGND.t345 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X384 a_5456_46# a_3177_n4294.t7 DGND.t402 DGND.t401 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X385 DGND.t24 A3.t6 a_2422_n1194# DGND.t23 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X386 DGND.t102 A7.t7 a_2422_n3674# DGND.t101 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X387 a_2422_n2068# B5.t7 a_2350_n2068# DVDD.t296 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X388 a_2995_n4294# a_2569_n4255# DGND.t63 DGND.t62 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X389 a_3226_n4062# a_2995_n4294# a_3368_n4255# DVDD.t46 sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X390 a_6023_n3054# A8.t6 DVDD.t28 DVDD.t27 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X391 DVDD.t179 B15.t7 a_4363_n828# DVDD.t178 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X392 a_143_n2276# a_2569_n1775# DGND.t125 DGND.t124 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X393 DVDD.t412 A12.t8 a_5855_n574# DVDD.t411 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X394 DGND.t424 A1.t6 a_2422_46# DGND.t423 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X395 DGND.t378 a_101_n1194# a_636_n1814# DGND.t377 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X396 DGND.t34 a_101_n3674# a_636_n4294# DGND.t33 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X397 a_6153_n2434# B8.t6 a_5402_n2306# DGND.t330 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X398 a_1557_46# B1.t5 a_1467_46# DGND.t193 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X399 a_185_n3674# a_143_n3516# a_101_n3674# DGND.t208 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X400 a_185_n1194# a_143_n1036# a_101_n1194# DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X401 a_101_46# B0.t7 a_11_412# DVDD.t404 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X402 a_5855_n1814# B14.t8 a_5773_n1814# DVDD.t53 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X403 DVDD.t143 a_636_n574# a_1997_412# DVDD.t142 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X404 a_143_n2276# a_2569_n1775# DVDD.t120 DVDD.t119 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X405 a_1201_n574# a_1261_n600# DGND.t190 DGND.t189 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X406 DVDD.t92 A7.t8 a_1291_n4294# DVDD.t91 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 a_4000_n2434# a_3946_n2306# a_3904_n2434# DGND.t322 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X408 DVDD.t374 a_101_n1194# a_636_n1814# DVDD.t373 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X409 a_3795_n2734# a_3765_n3080# a_3711_n2734# DGND.t523 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X410 DVDD.t219 a_143_n2276# a_541_n2068# DVDD.t218 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X411 a_1261_n600# A1.t7 DGND.t422 DGND.t421 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 a_185_n2434# B4.t6 DGND.t131 DGND.t130 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X413 a_1557_n2434# B5.t8 a_1467_n2068# DVDD.t19 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X414 a_1641_n2068# B5.t9 DVDD.t295 DVDD.t294 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X415 a_2908_n600# a_3874_n1220# a_3832_n1194# DGND.t133 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X416 a_3904_n3674# a_3874_n3700# a_3832_n3674# DGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X417 a_1997_n828# B3.t9 DVDD.t383 DVDD.t382 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X418 a_1291_n3054# a_1261_n3080# a_1201_n3054# DVDD.t222 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X419 a_4000_n2068# a_3874_n2460# DVDD.t260 DVDD.t259 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X420 a_3434_n4026# a_3946_n3546# DVDD.t264 DVDD.t263 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X421 a_1261_n3080# B5.t10 a_1647_n3054# DVDD.t289 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X422 a_2543_n2734# a_1201_n4294# a_2459_n2734# DGND.t461 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X423 a_894_412# Cin.t5 a_798_46# DVDD.t480 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X424 a_541_n3308# B6.t7 DVDD.t416 DVDD.t415 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X425 DGND.t140 a_636_n3054# a_1997_n2434# DGND.t139 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X426 a_101_n2434# B4.t7 a_11_n2434# DGND.t405 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X427 DVDD.t403 A9.t6 a_4697_n2068# DVDD.t402 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X428 DVDD.t445 a_n131_n1814# a_2273_n254# DVDD.t444 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X429 a_5402_n2306# a_2995_n4294# a_5819_n2434# DGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X430 a_2273_n2734# a_n131_n3054# DVDD.t469 DVDD.t468 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X431 a_798_46# a_101_46# a_541_412# DVDD.t80 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X432 a_2254_n3674# a_1557_n3674# a_1997_n3308# DVDD.t460 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X433 DGND.t38 A8.t7 a_5773_n3054# DGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X434 a_4691_n574# A13.t9 DVDD.t84 DVDD.t83 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X435 DVDD.t245 B13.t7 a_4363_412# DVDD.t244 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X436 DGND.t420 A1.t8 a_1641_46# DGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 a_5288_n3308# B10.t5 a_5192_n3308# DVDD.t246 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X438 a_1291_n4294# B7.t9 DVDD.t59 DVDD.t58 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X439 DVDD.t307 B8.t7 a_6023_n3054# DVDD.t306 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X440 a_1641_412# B1.t6 DVDD.t370 DVDD.t369 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X441 a_5288_46# B12.t6 a_5192_46# DGND.t404 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X442 DVDD.t156 B12.t7 a_5456_412# DVDD.t155 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X443 DVDD.t2 a_143_n1036# a_541_n828# DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X444 DGND.t240 A4.t6 a_185_n2434# DGND.t239 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X445 a_5819_n3674# A10.t7 DGND.t56 DGND.t55 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 a_5819_n1194# A14.t8 DGND.t348 DGND.t347 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X447 DVDD.t332 A9.t7 a_4000_n2068# DVDD.t331 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X448 a_2363_n254# a_n131_n574# a_2273_n254# DGND.t321 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X449 a_1647_n3054# A5.t7 DVDD.t372 DVDD.t371 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X450 a_5456_46# a_5402_174# a_5360_46# DGND.t349 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X451 a_2459_n2734# a_1201_n3054# a_2363_n2734# DGND.t501 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X452 a_6023_n4294# A10.t8 DVDD.t45 DVDD.t44 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 a_541_n3308# A6.t7 DVDD.t62 DVDD.t61 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X454 a_1479_n254# B1.t7 a_1201_n574# DGND.t475 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X455 DGND.t430 B8.t8 a_5456_n2434# DGND.t429 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X456 a_3736_n2434# A9.t8 DGND.t162 DGND.t161 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X457 DVDD.t439 B11.t9 a_4000_n3308# DVDD.t438 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X458 a_6153_n1194# B14.t9 a_5402_n1066# DGND.t329 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X459 a_6153_n3674# B10.t6 a_5402_n3546# DGND.t230 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 DGND.t20 A13.t10 a_4697_46# DGND.t19 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X461 a_3765_n600# B13.t8 a_4691_n254# DGND.t229 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X462 DVDD.t503 B10.t7 a_5819_n3308# DVDD.t502 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X463 a_3322_n4062# a_3861_n3080# a_3795_n2734# DGND.t203 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X464 DGND.t94 a_101_46# a_636_n574# DGND.t93 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X465 a_4523_n574# B13.t9 a_4441_n574# DVDD.t501 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X466 a_n71_n3080# A4.t7 DGND.t228 DGND.t227 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X467 a_315_n574# A0.t7 DVDD.t97 DVDD.t96 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X468 DGND.t122 B12.t8 a_5819_46# DGND.t121 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X469 a_4000_n1194# a_3946_n1066# a_2908_n600# DGND.t114 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X470 a_4000_n3674# a_3946_n3546# a_3904_n3674# DGND.t261 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X471 DVDD.t224 a_3669_n2822# a_3322_n4062# DVDD.t223 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X472 a_4441_n3054# B9.t9 DGND.t289 DGND.t288 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X473 DVDD.t422 A1.t9 a_1641_412# DVDD.t421 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X474 a_1467_n828# A3.t7 DVDD.t74 DVDD.t73 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X475 a_185_n1194# B2.t9 DGND.t127 DGND.t126 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X476 a_185_n3674# B6.t8 DGND.t411 DGND.t410 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X477 DVDD.t330 B14.t10 a_5819_n828# DVDD.t329 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X478 DVDD.t239 a_1557_46# a_143_n1036# DVDD.t238 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X479 DGND.t213 a_1557_n2434# a_143_n3516# DGND.t212 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X480 DGND.t181 A8.t8 a_6153_n2434# DGND.t180 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X481 a_5402_n1066# a_4204_n574# a_5819_n828# DVDD.t202 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X482 a_1291_n4294# a_1261_n4320# a_1201_n4294# DVDD.t376 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X483 a_3946_n1066# a_3874_n1220# a_4363_n828# DVDD.t126 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X484 a_1261_n4320# B7.t10 a_1647_n4294# DVDD.t60 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X485 a_2350_n3308# a_636_n4294# a_2254_n3674# DVDD.t22 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X486 a_5456_n2434# a_2995_n4294# DGND.t59 DGND.t58 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 a_541_n2068# B4.t8 DVDD.t158 DVDD.t157 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X488 DGND.t250 a_636_n1814# a_1997_n1194# DGND.t249 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X489 DGND.t29 a_636_n4294# a_1997_n3674# DGND.t28 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X490 a_101_n3674# B6.t9 a_11_n3674# DGND.t383 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X491 a_185_n828# B2.t10 DVDD.t118 DVDD.t117 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X492 a_3832_n828# B15.t8 a_3736_n828# DVDD.t393 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X493 a_101_n1194# B2.t11 a_11_n1194# DGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X494 a_5402_n1066# a_4204_n574# a_5819_n1194# DGND.t206 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X495 a_5402_n3546# a_4204_n3054# a_5819_n3674# DGND.t270 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 a_3368_n1775# a_3322_n1582# DVDD.t447 DVDD.t446 sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X497 a_5855_n3054# B8.t9 a_5773_n3054# DVDD.t93 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X498 a_2254_n2434# a_1557_n2434# a_1997_n2068# DVDD.t214 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X499 DGND.t67 A10.t9 a_5773_n4294# DGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X500 DGND.t396 A14.t9 a_5773_n1814# DGND.t395 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X501 a_5288_n2068# B8.t10 a_5192_n2068# DVDD.t72 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X502 a_5456_412# a_3177_n4294.t8 DVDD.t380 DVDD.t379 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X503 DVDD.t82 B10.t8 a_6023_n4294# DVDD.t81 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X504 DVDD.t315 a_101_n2434# a_636_n3054# DVDD.t314 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X505 a_3322_n4062# a_3543_n2822# DVDD.t509 DVDD.t508 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X506 a_798_n2434# a_101_n2434# a_541_n2434# DGND.t316 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X507 DGND.t392 A2.t6 a_185_n1194# DGND.t391 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X508 DGND.t226 A6.t8 a_185_n3674# DGND.t225 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 a_2543_n254# a_1201_n1814# a_2459_n254# DGND.t305 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 DGND.t83 A13.t11 a_4441_n574# DGND.t82 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X511 a_1557_n1194# B3.t10 a_1467_n828# DVDD.t165 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X512 DVDD.t392 A14.t10 a_5855_n1814# DVDD.t391 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X513 DGND.t87 B0.t8 a_n71_n600# DGND.t86 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X514 a_4204_n574# a_3946_174# DVDD.t351 DVDD.t350 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X515 a_5456_n3308# a_5402_n3546# a_5360_n3674# DVDD.t241 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X516 a_1647_n4294# A7.t9 DVDD.t88 DVDD.t87 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 DGND.t147 a_4441_n574# a_3765_n600# DGND.t146 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X518 a_3832_n2434# B9.t10 a_3736_n2434# DGND.t510 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X519 a_1997_n2434# B5.t11 DGND.t129 DGND.t128 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X520 DVDD.t301 a_n131_n4294# a_2273_n2734# DVDD.t300 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X521 DVDD.t90 A7.t10 a_2422_n3308# DVDD.t89 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X522 a_3368_n4255# a_3322_n4062# DVDD.t191 DVDD.t190 sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X523 a_3946_n2306# a_3874_n2460# a_4363_n2434# DGND.t257 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X524 a_541_n2068# A4.t8 DVDD.t500 DVDD.t499 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 a_541_46# A0.t8 DGND.t447 DGND.t446 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X526 DGND.t247 B14.t11 a_5456_n1194# DGND.t246 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X527 a_3736_n3674# A11.t10 DGND.t277 DGND.t276 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X528 DGND.t18 B10.t9 a_5456_n3674# DGND.t17 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X529 a_3736_n1194# A15.t9 DGND.t51 DGND.t50 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X530 a_3368_n3928# a_3322_n4062# DGND.t197 DGND.t196 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X531 a_3368_n1448# a_3322_n1582# DGND.t455 DGND.t454 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X532 a_5456_n828# a_4204_n574# DVDD.t201 DVDD.t200 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X533 DVDD.t513 B9.t11 a_4000_n2068# DVDD.t512 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X534 DGND.t375 A12.t9 a_6153_46# DGND.t374 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X535 a_3861_n600# B12.t9 a_6023_n254# DGND.t11 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X536 a_185_n3308# a_143_n3516# a_101_n3674# DVDD.t210 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X537 DVDD.t234 B8.t11 a_5819_n2068# DVDD.t233 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X538 a_185_n828# a_143_n1036# a_101_n1194# DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 a_1997_n2434# A5.t8 DGND.t479 DGND.t478 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X540 DGND.t520 B13.t10 a_4363_46# DGND.t519 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X541 DGND.t304 a_2908_n600# S15.t0 DGND.t303 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X542 a_n71_n1840# A2.t7 DGND.t394 DGND.t393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X543 a_n71_n4320# A6.t9 DGND.t77 DGND.t76 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X544 DGND.t518 A4.t9 a_966_n2434# DGND.t517 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X545 a_2422_412# B1.t8 a_2350_412# DVDD.t291 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X546 a_3589_n3928# a_2995_n4294# a_3226_n4062# DGND.t57 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X547 a_4441_n4294# B11.t10 DGND.t451 DGND.t450 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X548 a_4441_n1814# B15.t9 DGND.t432 DGND.t431 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X549 a_3589_n1448# a_3177_n4294.t9 a_3226_n1582# DGND.t47 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X550 DGND.t353 A14.t11 a_6153_n1194# DGND.t352 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X551 DGND.t398 a_1557_n1194# a_1968_n1814# DGND.t397 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X552 DGND.t69 A10.t10 a_6153_n3674# DGND.t68 sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X553 DGND.t470 a_1557_n3674# a_1968_n4294# DGND.t469 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X554 a_3904_n3674# a_3874_n3700# a_3832_n3308# DVDD.t484 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X555 a_4363_n2434# A9.t9 DGND.t500 DGND.t499 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X556 DGND.t522 A4.t10 a_147_n2734# DGND.t521 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X557 a_541_412# A0.t9 DVDD.t431 DVDD.t430 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X558 a_5456_n1194# a_4204_n574# DGND.t205 DGND.t204 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X559 a_5456_n3674# a_4204_n3054# DGND.t269 DGND.t268 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X560 a_2350_n2068# a_636_n3054# a_2254_n2434# DVDD.t130 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X561 a_315_n1814# A2.t8 DVDD.t185 DVDD.t184 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X562 a_3711_n254# a_3669_n342# a_3627_n254# DGND.t248 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X563 a_185_46# Cin.t6 a_101_46# DGND.t179 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X564 DGND.t46 A0.t10 a_147_n254# DGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X565 a_4691_n2734# A9.t10 DGND.t369 DGND.t368 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X566 a_4523_n1814# B15.t10 a_4441_n1814# DVDD.t237 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X567 DVDD.t420 A1.t10 a_2422_412# DVDD.t419 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X568 a_1647_n574# A1.t11 DVDD.t418 DVDD.t417 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X569 a_3669_n342# a_4441_n1814# a_4691_n1814# DVDD.t136 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X570 a_5855_n4294# B10.t10 a_5773_n4294# DVDD.t67 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X571 a_1997_n828# A3.t8 DVDD.t152 DVDD.t151 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X572 DVDD.t397 a_1557_n1194# a_1968_n1814# DVDD.t396 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X573 a_5819_412# A12.t10 DVDD.t161 DVDD.t160 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X574 a_2995_n4294# a_2569_n4255# DVDD.t52 DVDD.t51 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X575 DGND.t409 A8.t9 a_5456_n2434# DGND.t408 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X576 a_894_n2434# a_143_n2276# a_798_n2434# DGND.t215 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X577 a_1291_n574# a_1261_n600# a_1201_n574# DVDD.t186 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X578 DVDD.t337 A3.t9 a_2422_n828# DVDD.t336 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X579 a_1641_46# B1.t9 DGND.t413 DGND.t412 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X580 DVDD.t25 a_101_n3674# a_636_n4294# DVDD.t24 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X581 a_3685_n1775# a_3434_n1546# a_3226_n1582# DVDD.t297 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X582 a_185_46# B0.t9 DGND.t42 DGND.t41 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X583 a_3946_174# a_3874_20# a_4363_46# DGND.t264 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X584 a_798_n1194# a_101_n1194# a_541_n1194# DGND.t376 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X585 a_798_n3674# a_101_n3674# a_541_n3674# DGND.t32 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X586 DVDD.t355 a_2273_n254# a_2315_n1775# DVDD.t354 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X587 a_3874_n2460# a_5402_n2306# DGND.t201 DGND.t200 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X588 a_11_n2434# A4.t11 DGND.t534 DGND.t533 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X589 a_5819_n3308# A10.t11 DVDD.t516 DVDD.t515 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X590 a_11_412# A0.t11 DVDD.t95 DVDD.t94 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X591 a_101_46# B0.t10 a_11_46# DGND.t336 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X592 a_4000_n828# a_3874_n1220# DVDD.t125 DVDD.t124 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X593 a_147_n2734# B4.t9 a_n131_n3054# DGND.t298 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X594 a_5456_n2068# a_5402_n2306# a_5360_n2434# DVDD.t194 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X595 a_1997_n1194# B3.t11 DGND.t15 DGND.t14 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X596 a_3832_n1194# B15.t11 a_3736_n1194# DGND.t92 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X597 a_3832_n3674# B11.t11 a_3736_n3674# DGND.t443 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X598 a_1997_n3674# B7.t11 DGND.t245 DGND.t244 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X599 DGND.t309 B4.t10 a_n71_n3080# DGND.t308 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X600 a_3226_n4062# a_3434_n4026# a_3368_n3928# DGND.t158 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X601 a_3226_n1582# a_3434_n1546# a_3368_n1448# DGND.t295 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X602 a_5456_n828# a_5402_n1066# a_5360_n1194# DVDD.t528 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X603 DVDD.t55 A5.t9 a_2422_n2068# DVDD.t54 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X604 a_3946_n1066# a_3874_n1220# a_4363_n1194# DGND.t132 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X605 a_3946_n3546# a_3874_n3700# a_4363_n3674# DGND.t481 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X606 a_3322_n4062# a_3765_n3080# DVDD.t527 DVDD.t526 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X607 a_966_n2434# B4.t11 a_894_n2434# DGND.t123 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X608 DGND.t360 A9.t11 a_4441_n3054# DGND.t359 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X609 a_4000_n828# a_3946_n1066# a_2908_n600# DVDD.t110 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X610 a_5192_n2434# A8.t10 DGND.t104 DGND.t103 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X611 DVDD.t511 a_3655_n1516# a_3685_n1775# DVDD.t510 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X612 DVDD.t498 Cin.t7 a_541_412# DVDD.t497 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X613 a_2273_n254# a_n131_n574# DVDD.t320 DVDD.t319 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X614 a_6153_n3308# B10.t11 a_5402_n3546# DVDD.t335 sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X615 DGND.t371 A5.t10 a_1641_n2434# DGND.t370 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X616 a_2273_n2734# a_1201_n4294# DVDD.t456 DVDD.t455 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X617 a_3685_n4255# a_3434_n4026# a_3226_n4062# DVDD.t162 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X618 a_185_n2068# a_143_n2276# a_101_n2434# DVDD.t217 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X619 a_1997_n1194# A3.t10 DGND.t332 DGND.t331 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 a_1997_n3674# A7.t11 DGND.t89 DGND.t88 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X621 DVDD.t147 a_2273_n2734# a_2315_n4255# DVDD.t146 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X622 a_1291_n574# B1.t10 DVDD.t362 DVDD.t361 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X623 DGND.t224 a_3655_n3996# a_3589_n3928# DGND.t223 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X624 DGND.t507 a_3655_n1516# a_3589_n1448# DGND.t506 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X625 a_1997_412# B1.t11 DVDD.t478 DVDD.t477 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X626 DVDD.t17 B12.t10 a_5819_412# DVDD.t16 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X627 DGND.t326 a_3226_n4062# a_3177_n4294.t0 DGND.t325 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X628 DVDD.t167 A8.t11 a_5855_n3054# DVDD.t166 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 DGND.t382 a_3226_n1582# a_3177_n1814# DGND.t381 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X630 DGND.t362 a_2273_n254# a_2315_n1775# DGND.t361 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X631 DGND.t153 a_2273_n2734# a_2315_n4255# DGND.t152 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X632 DVDD.t177 A3.t11 a_1641_n828# DVDD.t176 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X633 DGND.t188 A2.t9 a_966_n1194# DGND.t187 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X634 DGND.t75 A6.t10 a_966_n3674# DGND.t74 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X635 a_4000_n3308# a_3946_n3546# a_3904_n3674# DVDD.t262 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X636 a_4000_412# a_3946_174# a_3904_46# DVDD.t349 sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X637 a_185_412# B0.t11 DVDD.t69 DVDD.t68 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X638 a_5819_46# A12.t11 DGND.t313 DGND.t312 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X639 a_185_n3308# B6.t10 DVDD.t366 DVDD.t365 sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X640 a_5773_n574# B12.t11 DGND.t157 DGND.t156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X641 a_2350_n828# a_636_n1814# a_2254_n1194# DVDD.t251 sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X642 a_3736_n828# A15.t10 DVDD.t41 DVDD.t40 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X643 DVDD.t518 B13.t11 a_4691_n574# DVDD.t517 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X644 a_4363_n1194# A15.t11 DGND.t177 DGND.t176 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X645 a_4363_n3674# A11.t11 DGND.t275 DGND.t274 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X646 a_3904_n2434# a_3874_n2460# a_3832_n2068# DVDD.t258 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X647 a_3904_46# a_3874_20# a_3832_412# DVDD.t265 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X648 a_3322_n1582# a_3861_n600# a_3795_n254# DGND.t458 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X649 DGND.t49 A2.t10 a_147_n1494# DGND.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X650 DGND.t165 A6.t11 a_147_n3974# DGND.t164 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X651 a_1467_n2434# A5.t11 DGND.t498 DGND.t497 sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X652 DVDD.t39 A2.t11 a_966_n828# DVDD.t38 sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X653 DVDD.t79 a_101_46# a_636_n574# DVDD.t78 sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X654 DVDD.t231 a_3655_n3996# a_3685_n4255# DVDD.t230 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X655 DVDD.t378 a_3226_n1582# a_3177_n1814# DVDD.t377 sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X656 DVDD.t21 a_636_n4294# a_1997_n3308# DVDD.t20 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X657 a_101_n3674# B6.t11 a_11_n3308# DVDD.t13 sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
R0 A11.n2 A11.t9 373.283
R1 A11.n1 A11.t2 347.577
R2 A11.n0 A11.t8 334.723
R3 A11.n4 A11.t3 323.476
R4 A11.n4 A11.t11 217.436
R5 A11.n6 A11.t5 212.081
R6 A11.n7 A11.t7 212.081
R7 A11.n0 A11.t4 206.19
R8 A11.n1 A11.t10 193.337
R9 A11.n9 A11.n8 174.552
R10 A11.n5 A11.n4 169.833
R11 A11.n2 A11.t6 167.63
R12 A11.n3 A11.n1 166.843
R13 A11.n3 A11.n2 166.421
R14 A11.n10 A11.n0 152
R15 A11.n6 A11.t0 139.78
R16 A11.n7 A11.t1 139.78
R17 A11.n8 A11.n6 37.246
R18 A11.n8 A11.n7 24.1005
R19 A11.n10 A11.n9 17.5294
R20 A11.n10 A11 14.0805
R21 A11 A11.n10 2.51479
R22 A11.n5 A11.n3 1.55989
R23 A11.n9 A11.n5 0.112749
R24 DGND.n811 DGND.n810 8899.17
R25 DGND.n433 DGND.t303 3347.83
R26 DGND.t124 DGND.t381 1942.47
R27 DGND.t136 DGND.n433 1721.74
R28 DGND.t452 DGND.n951 1721.74
R29 DGND.t517 DGND.t220 1714.38
R30 DGND.t272 DGND.t365 1714.38
R31 DGND.t74 DGND.t379 1714.38
R32 DGND.t487 DGND.t103 1714.38
R33 DGND.t495 DGND.t144 1714.38
R34 DGND.t427 DGND.t187 1714.38
R35 DGND.t169 DGND.t146 1714.38
R36 DGND.t286 DGND.t189 1714.38
R37 DGND.n810 DGND.n203 1444.51
R38 DGND.t296 DGND.t128 1383.28
R39 DGND.t463 DGND.t459 1383.28
R40 DGND.t293 DGND.t244 1383.28
R41 DGND.t327 DGND.t540 1383.28
R42 DGND.t119 DGND.t333 1383.28
R43 DGND.t14 DGND.t508 1383.28
R44 DGND.t519 DGND.t191 1383.28
R45 DGND.t412 DGND.t291 1383.28
R46 DGND.t220 DGND.t497 1265.55
R47 DGND.t365 DGND.t280 1265.55
R48 DGND.t379 DGND.t385 1265.55
R49 DGND.t98 DGND.t487 1265.55
R50 DGND.t144 DGND.t476 1265.55
R51 DGND.t112 DGND.t427 1265.55
R52 DGND.t146 DGND.t19 1265.55
R53 DGND.t189 DGND.t414 1265.55
R54 DGND.n433 DGND.n432 1215.29
R55 DGND.n156 DGND.n155 1202
R56 DGND.n892 DGND.n891 1202
R57 DGND.n813 DGND.n812 1202
R58 DGND.n894 DGND.n893 1202
R59 DGND.n316 DGND.n315 1202
R60 DGND.n809 DGND.n808 1202
R61 DGND.n608 DGND.n607 1202
R62 DGND.n688 DGND.n687 1202
R63 DGND.n606 DGND.n605 1202
R64 DGND.n690 DGND.n689 1202
R65 DGND.n951 DGND.n950 1202
R66 DGND.n953 DGND.n952 1202
R67 DGND.n435 DGND.n434 1202
R68 DGND.t310 DGND.t308 1044.82
R69 DGND.t17 DGND.t231 1044.82
R70 DGND.t117 DGND.t182 1044.82
R71 DGND.t429 DGND.t90 1044.82
R72 DGND.t246 DGND.t64 1044.82
R73 DGND.t441 DGND.t9 1044.82
R74 DGND.t242 DGND.t156 1044.82
R75 DGND.t167 DGND.t86 1044.82
R76 DGND.n810 DGND.t301 971.237
R77 DGND.t325 DGND.n811 971.237
R78 DGND.n811 DGND.t62 971.237
R79 DGND.n810 DGND.t504 971.237
R80 DGND.t57 DGND.t158 919.732
R81 DGND.t217 DGND.t466 919.732
R82 DGND.t47 DGND.t295 919.732
R83 DGND.t54 DGND.t341 919.732
R84 DGND.t196 DGND.t325 802.008
R85 DGND.t62 DGND.t154 802.008
R86 DGND.t381 DGND.t454 802.008
R87 DGND.t363 DGND.t124 802.008
R88 DGND.t214 DGND.t141 706.355
R89 DGND.t215 DGND.t316 706.355
R90 DGND.t271 DGND.t236 706.355
R91 DGND.t261 DGND.t482 706.355
R92 DGND.t443 DGND.t276 706.355
R93 DGND.t223 DGND.t57 706.355
R94 DGND.t4 DGND.t217 706.355
R95 DGND.t335 DGND.t101 706.355
R96 DGND.t471 DGND.t30 706.355
R97 DGND.t211 DGND.t32 706.355
R98 DGND.t61 DGND.t202 706.355
R99 DGND.t258 DGND.t322 706.355
R100 DGND.t207 DGND.t524 706.355
R101 DGND.t114 DGND.t133 706.355
R102 DGND.t92 DGND.t50 706.355
R103 DGND.t506 DGND.t47 706.355
R104 DGND.t341 DGND.t357 706.355
R105 DGND.t23 DGND.t241 706.355
R106 DGND.t251 DGND.t399 706.355
R107 DGND.t3 DGND.t376 706.355
R108 DGND.t511 DGND.t349 706.355
R109 DGND.t356 DGND.t265 706.355
R110 DGND.t235 DGND.t151 706.355
R111 DGND.t403 DGND.t95 706.355
R112 DGND.t405 DGND.t533 662.207
R113 DGND.t230 DGND.t68 662.207
R114 DGND.t383 DGND.t35 662.207
R115 DGND.t330 DGND.t180 662.207
R116 DGND.t329 DGND.t352 662.207
R117 DGND.t8 DGND.t467 662.207
R118 DGND.t290 DGND.t374 662.207
R119 DGND.t336 DGND.t71 662.207
R120 DGND.t478 DGND.t214 654.85
R121 DGND.t278 DGND.t261 654.85
R122 DGND.t88 DGND.t471 654.85
R123 DGND.t322 DGND.t515 654.85
R124 DGND.t253 DGND.t114 654.85
R125 DGND.t399 DGND.t331 654.85
R126 DGND.t433 DGND.t356 654.85
R127 DGND.t444 DGND.t235 654.85
R128 DGND.t461 DGND.t301 618.061
R129 DGND.t139 DGND.t478 618.061
R130 DGND.t535 DGND.t218 618.061
R131 DGND.t218 DGND.t310 618.061
R132 DGND.t268 DGND.t17 618.061
R133 DGND.t159 DGND.t268 618.061
R134 DGND.t483 DGND.t278 618.061
R135 DGND.t28 DGND.t88 618.061
R136 DGND.t194 DGND.t209 618.061
R137 DGND.t209 DGND.t117 618.061
R138 DGND.t58 DGND.t429 618.061
R139 DGND.t408 DGND.t58 618.061
R140 DGND.t515 DGND.t259 618.061
R141 DGND.t504 DGND.t222 618.061
R142 DGND.t204 DGND.t246 618.061
R143 DGND.t339 DGND.t204 618.061
R144 DGND.t134 DGND.t253 618.061
R145 DGND.t331 DGND.t249 618.061
R146 DGND.t319 DGND.t1 618.061
R147 DGND.t1 DGND.t441 618.061
R148 DGND.t401 DGND.t242 618.061
R149 DGND.t26 DGND.t401 618.061
R150 DGND.t266 DGND.t433 618.061
R151 DGND.t248 DGND.t136 618.061
R152 DGND.t305 DGND.t452 618.061
R153 DGND.t149 DGND.t444 618.061
R154 DGND.t446 DGND.t345 618.061
R155 DGND.t345 DGND.t167 618.061
R156 DGND.t316 DGND.t317 588.63
R157 DGND.t236 DGND.t237 588.63
R158 DGND.t32 DGND.t33 588.63
R159 DGND.t202 DGND.t200 588.63
R160 DGND.t524 DGND.t525 588.63
R161 DGND.t376 DGND.t377 588.63
R162 DGND.t349 DGND.t350 588.63
R163 DGND.t95 DGND.t93 588.63
R164 DGND.t417 DGND.t296 573.913
R165 DGND.t337 DGND.t370 573.913
R166 DGND.t372 DGND.t142 573.913
R167 DGND.t306 DGND.t186 573.913
R168 DGND.t462 DGND.t465 573.913
R169 DGND.t284 DGND.t481 573.913
R170 DGND.t282 DGND.t274 573.913
R171 DGND.t450 DGND.t463 573.913
R172 DGND.t513 DGND.t293 573.913
R173 DGND.t43 DGND.t184 573.913
R174 DGND.t387 DGND.t31 573.913
R175 DGND.t175 DGND.t367 573.913
R176 DGND.t344 DGND.t512 573.913
R177 DGND.t257 DGND.t368 573.913
R178 DGND.t499 DGND.t359 573.913
R179 DGND.t540 DGND.t288 573.913
R180 DGND.t25 DGND.t97 573.913
R181 DGND.t389 DGND.t132 573.913
R182 DGND.t342 DGND.t176 573.913
R183 DGND.t431 DGND.t119 573.913
R184 DGND.t508 DGND.t6 573.913
R185 DGND.t439 DGND.t502 573.913
R186 DGND.t252 DGND.t437 573.913
R187 DGND.t384 DGND.t73 573.913
R188 DGND.t229 DGND.t480 573.913
R189 DGND.t435 DGND.t264 573.913
R190 DGND.t82 DGND.t39 573.913
R191 DGND.t537 DGND.t519 573.913
R192 DGND.t108 DGND.t412 573.913
R193 DGND.t421 DGND.t419 573.913
R194 DGND.t425 DGND.t148 573.913
R195 DGND.t475 DGND.t193 573.913
R196 DGND.n951 DGND.t303 566.556
R197 DGND.t123 DGND.t215 529.766
R198 DGND.t100 DGND.t271 529.766
R199 DGND.t472 DGND.t211 529.766
R200 DGND.t539 DGND.t61 529.766
R201 DGND.t529 DGND.t207 529.766
R202 DGND.t416 DGND.t3 529.766
R203 DGND.t404 DGND.t511 529.766
R204 DGND.t138 DGND.t403 529.766
R205 DGND.n812 DGND.t158 522.409
R206 DGND.t466 DGND.n892 522.409
R207 DGND.t295 DGND.n688 522.409
R208 DGND.n607 DGND.t54 522.409
R209 DGND.t501 DGND.t531 434.115
R210 DGND.t474 DGND.t307 434.115
R211 DGND.t510 DGND.t203 434.115
R212 DGND.t161 DGND.t523 434.115
R213 DGND.t458 DGND.t473 434.115
R214 DGND.t400 DGND.t84 434.115
R215 DGND.t143 DGND.t423 434.115
R216 DGND.t321 DGND.t163 434.115
R217 DGND.n155 DGND.t123 404.683
R218 DGND.n315 DGND.t100 404.683
R219 DGND.n893 DGND.t472 404.683
R220 DGND.n809 DGND.t539 404.683
R221 DGND.n689 DGND.t529 404.683
R222 DGND.n606 DGND.t416 404.683
R223 DGND.n434 DGND.t404 404.683
R224 DGND.n952 DGND.t138 404.683
R225 DGND.t128 DGND.t212 389.967
R226 DGND.t459 DGND.t262 389.967
R227 DGND.t244 DGND.t469 389.967
R228 DGND.t323 DGND.t327 389.967
R229 DGND.t333 DGND.t115 389.967
R230 DGND.t397 DGND.t14 389.967
R231 DGND.t191 DGND.t354 389.967
R232 DGND.t291 DGND.t233 389.967
R233 DGND.t482 DGND.t198 375.252
R234 DGND.t276 DGND.t223 375.252
R235 DGND.t101 DGND.t4 375.252
R236 DGND.t30 DGND.t152 375.252
R237 DGND.t133 DGND.t456 375.252
R238 DGND.t50 DGND.t506 375.252
R239 DGND.t357 DGND.t23 375.252
R240 DGND.t361 DGND.t251 375.252
R241 DGND.t533 DGND.t314 353.178
R242 DGND.t68 DGND.t255 353.178
R243 DGND.t35 DGND.t489 353.178
R244 DGND.t180 DGND.t406 353.178
R245 DGND.t352 DGND.t171 353.178
R246 DGND.t467 DGND.t52 353.178
R247 DGND.t374 DGND.t173 353.178
R248 DGND.t71 DGND.t527 353.178
R249 DGND.t308 DGND.t130 338.462
R250 DGND.t227 DGND.t239 338.462
R251 DGND.t521 DGND.t216 338.462
R252 DGND.t298 DGND.t405 338.462
R253 DGND.t105 DGND.t230 338.462
R254 DGND.t106 DGND.t270 338.462
R255 DGND.t66 DGND.t55 338.462
R256 DGND.t231 DGND.t80 338.462
R257 DGND.t182 DGND.t410 338.462
R258 DGND.t76 DGND.t225 338.462
R259 DGND.t164 DGND.t208 338.462
R260 DGND.t178 DGND.t383 338.462
R261 DGND.t96 DGND.t330 338.462
R262 DGND.t78 DGND.t60 338.462
R263 DGND.t37 DGND.t110 338.462
R264 DGND.t90 DGND.t21 338.462
R265 DGND.t530 DGND.t329 338.462
R266 DGND.t491 DGND.t206 338.462
R267 DGND.t395 DGND.t347 338.462
R268 DGND.t64 DGND.t485 338.462
R269 DGND.t9 DGND.t126 338.462
R270 DGND.t393 DGND.t391 338.462
R271 DGND.t48 DGND.t0 338.462
R272 DGND.t16 DGND.t8 338.462
R273 DGND.t11 DGND.t290 338.462
R274 DGND.t12 DGND.t70 338.462
R275 DGND.t299 DGND.t312 338.462
R276 DGND.t156 DGND.t121 338.462
R277 DGND.t86 DGND.t41 338.462
R278 DGND.t448 DGND.t493 338.462
R279 DGND.t45 DGND.t179 338.462
R280 DGND.t166 DGND.t336 338.462
R281 DGND.n155 DGND.t517 301.673
R282 DGND.n315 DGND.t272 301.673
R283 DGND.n893 DGND.t74 301.673
R284 DGND.t103 DGND.n809 301.673
R285 DGND.n689 DGND.t495 301.673
R286 DGND.t187 DGND.n606 301.673
R287 DGND.n434 DGND.t169 301.673
R288 DGND.n952 DGND.t286 301.673
R289 DGND.t130 DGND.t227 279.599
R290 DGND.t239 DGND.t521 279.599
R291 DGND.t216 DGND.t298 279.599
R292 DGND.t270 DGND.t105 279.599
R293 DGND.t55 DGND.t106 279.599
R294 DGND.t80 DGND.t66 279.599
R295 DGND.t410 DGND.t76 279.599
R296 DGND.t225 DGND.t164 279.599
R297 DGND.t208 DGND.t178 279.599
R298 DGND.t60 DGND.t96 279.599
R299 DGND.t110 DGND.t78 279.599
R300 DGND.t21 DGND.t37 279.599
R301 DGND.t206 DGND.t530 279.599
R302 DGND.t347 DGND.t491 279.599
R303 DGND.t485 DGND.t395 279.599
R304 DGND.t126 DGND.t393 279.599
R305 DGND.t391 DGND.t48 279.599
R306 DGND.t0 DGND.t16 279.599
R307 DGND.t70 DGND.t11 279.599
R308 DGND.t312 DGND.t12 279.599
R309 DGND.t121 DGND.t299 279.599
R310 DGND.t41 DGND.t448 279.599
R311 DGND.t493 DGND.t45 279.599
R312 DGND.t179 DGND.t166 279.599
R313 DGND.n52 DGND.t183 278.589
R314 DGND.n842 DGND.t514 278.589
R315 DGND.n214 DGND.t451 278.589
R316 DGND.n297 DGND.t232 278.589
R317 DGND.n123 DGND.t309 278.589
R318 DGND.n106 DGND.t418 278.589
R319 DGND.n749 DGND.t289 278.589
R320 DGND.n705 DGND.t91 278.589
R321 DGND.n572 DGND.t10 278.589
R322 DGND.n500 DGND.t7 278.589
R323 DGND.n649 DGND.t432 278.589
R324 DGND.n468 DGND.t65 278.589
R325 DGND.n6 DGND.t87 278.589
R326 DGND.n33 DGND.t109 278.589
R327 DGND.n397 DGND.t538 278.589
R328 DGND.n349 DGND.t157 278.589
R329 DGND.t307 DGND.t501 272.241
R330 DGND.t523 DGND.t510 272.241
R331 DGND.t473 DGND.t400 272.241
R332 DGND.t163 DGND.t143 272.241
R333 DGND.n62 DGND.t36 259.74
R334 DGND.n845 DGND.t386 259.74
R335 DGND.n211 DGND.t281 259.74
R336 DGND.n285 DGND.t69 259.74
R337 DGND.n133 DGND.t534 259.74
R338 DGND.n109 DGND.t498 259.74
R339 DGND.n746 DGND.t99 259.74
R340 DGND.n714 DGND.t181 259.74
R341 DGND.n582 DGND.t468 259.74
R342 DGND.n553 DGND.t113 259.74
R343 DGND.n634 DGND.t477 259.74
R344 DGND.n456 DGND.t353 259.74
R345 DGND.n980 DGND.t72 259.74
R346 DGND.n36 DGND.t415 259.74
R347 DGND.n389 DGND.t20 259.74
R348 DGND.n337 DGND.t375 259.74
R349 DGND.n73 DGND.t118 239.281
R350 DGND.n835 DGND.t245 239.281
R351 DGND.n221 DGND.t460 239.281
R352 DGND.n302 DGND.t18 239.281
R353 DGND.n144 DGND.t311 239.281
R354 DGND.n99 DGND.t129 239.281
R355 DGND.n756 DGND.t328 239.281
R356 DGND.n703 DGND.t430 239.281
R357 DGND.n593 DGND.t442 239.281
R358 DGND.n531 DGND.t15 239.281
R359 DGND.n654 DGND.t334 239.281
R360 DGND.n473 DGND.t247 239.281
R361 DGND.n965 DGND.t168 239.281
R362 DGND.n26 DGND.t292 239.281
R363 DGND.n404 DGND.t192 239.281
R364 DGND.n354 DGND.t243 239.281
R365 DGND.n898 DGND.t75 237.536
R366 DGND.n883 DGND.t102 237.536
R367 DGND.n239 DGND.t277 237.536
R368 DGND.n320 DGND.t273 237.536
R369 DGND.n160 DGND.t518 237.536
R370 DGND.n197 DGND.t532 237.536
R371 DGND.n770 DGND.t162 237.536
R372 DGND.n805 DGND.t104 237.536
R373 DGND.n562 DGND.t188 237.536
R374 DGND.n520 DGND.t24 237.536
R375 DGND.n678 DGND.t51 237.536
R376 DGND.n694 DGND.t496 237.536
R377 DGND.n906 DGND.t287 237.536
R378 DGND.n943 DGND.t424 237.536
R379 DGND.n422 DGND.t85 237.536
R380 DGND.n439 DGND.t170 237.536
R381 DGND.t212 DGND.t139 228.095
R382 DGND.t262 DGND.t483 228.095
R383 DGND.t469 DGND.t28 228.095
R384 DGND.t259 DGND.t323 228.095
R385 DGND.t115 DGND.t134 228.095
R386 DGND.t249 DGND.t397 228.095
R387 DGND.t354 DGND.t266 228.095
R388 DGND.t233 DGND.t149 228.095
R389 DGND.n55 DGND.n54 200.127
R390 DGND.n859 DGND.n858 200.127
R391 DGND.n262 DGND.n261 200.127
R392 DGND.n296 DGND.n282 200.127
R393 DGND.n126 DGND.n125 200.127
R394 DGND.n173 DGND.n172 200.127
R395 DGND.n793 DGND.n792 200.127
R396 DGND.n720 DGND.n709 200.127
R397 DGND.n575 DGND.n574 200.127
R398 DGND.n547 DGND.n499 200.127
R399 DGND.n627 DGND.n626 200.127
R400 DGND.n467 DGND.n453 200.127
R401 DGND.n973 DGND.n5 200.127
R402 DGND.n919 DGND.n918 200.127
R403 DGND.n395 DGND.n381 200.127
R404 DGND.n348 DGND.n334 200.127
R405 DGND.n821 DGND.n820 199.739
R406 DGND.n817 DGND.n88 199.739
R407 DGND.n613 DGND.n612 199.739
R408 DGND.n684 DGND.n615 199.739
R409 DGND.n46 DGND.n45 198.964
R410 DGND.n51 DGND.n50 198.964
R411 DGND.n874 DGND.n833 198.964
R412 DGND.n864 DGND.n838 198.964
R413 DGND.n256 DGND.n216 198.964
R414 DGND.n248 DGND.n223 198.964
R415 DGND.n280 DGND.n279 198.964
R416 DGND.n276 DGND.n275 198.964
R417 DGND.n117 DGND.n116 198.964
R418 DGND.n122 DGND.n121 198.964
R419 DGND.n188 DGND.n97 198.964
R420 DGND.n178 DGND.n102 198.964
R421 DGND.n787 DGND.n751 198.964
R422 DGND.n779 DGND.n758 198.964
R423 DGND.n724 DGND.n723 198.964
R424 DGND.n732 DGND.n730 198.964
R425 DGND.n565 DGND.n564 198.964
R426 DGND.n571 DGND.n570 198.964
R427 DGND.n533 DGND.n530 198.964
R428 DGND.n542 DGND.n541 198.964
R429 DGND.n643 DGND.n642 198.964
R430 DGND.n656 DGND.n655 198.964
R431 DGND.n451 DGND.n450 198.964
R432 DGND.n447 DGND.n446 198.964
R433 DGND.n9 DGND.n8 198.964
R434 DGND.n969 DGND.n967 198.964
R435 DGND.n934 DGND.n24 198.964
R436 DGND.n924 DGND.n29 198.964
R437 DGND.n402 DGND.n401 198.964
R438 DGND.n413 DGND.n374 198.964
R439 DGND.n332 DGND.n331 198.964
R440 DGND.n328 DGND.n327 198.964
R441 DGND.n831 DGND.n830 185
R442 DGND.n829 DGND.n823 185
R443 DGND.n234 DGND.n233 185
R444 DGND.n232 DGND.n226 185
R445 DGND.n514 DGND.n508 185
R446 DGND.n516 DGND.n515 185
R447 DGND.n674 DGND.n673 185
R448 DGND.n672 DGND.n670 185
R449 DGND.t531 DGND.t461 183.946
R450 DGND.n812 DGND.t196 183.946
R451 DGND.n892 DGND.t154 183.946
R452 DGND.t222 DGND.t161 183.946
R453 DGND.n688 DGND.t454 183.946
R454 DGND.n607 DGND.t363 183.946
R455 DGND.t84 DGND.t248 183.946
R456 DGND.t423 DGND.t305 183.946
R457 DGND.n48 DGND.t34 158.361
R458 DGND.n869 DGND.t470 158.361
R459 DGND.n219 DGND.t263 158.361
R460 DGND.n306 DGND.t238 158.361
R461 DGND.n119 DGND.t318 158.361
R462 DGND.n183 DGND.t213 158.361
R463 DGND.n754 DGND.t324 158.361
R464 DGND.n736 DGND.t201 158.361
R465 DGND.n568 DGND.t378 158.361
R466 DGND.n504 DGND.t398 158.361
R467 DGND.n661 DGND.t116 158.361
R468 DGND.n477 DGND.t526 158.361
R469 DGND.n11 DGND.t94 158.361
R470 DGND.n929 DGND.t234 158.361
R471 DGND.n430 DGND.t304 158.361
R472 DGND.n410 DGND.t355 158.361
R473 DGND.n358 DGND.t351 158.361
R474 DGND.t198 DGND.t443 154.516
R475 DGND.t152 DGND.t335 154.516
R476 DGND.t456 DGND.t92 154.516
R477 DGND.t241 DGND.t361 154.516
R478 DGND.n201 DGND.t302 149.493
R479 DGND.n767 DGND.t505 149.493
R480 DGND.n947 DGND.t453 149.493
R481 DGND.n426 DGND.t137 149.493
R482 DGND.n61 DGND.t490 144.886
R483 DGND.n847 DGND.t380 144.886
R484 DGND.n271 DGND.t366 144.886
R485 DGND.n287 DGND.t256 144.886
R486 DGND.n132 DGND.t315 144.886
R487 DGND.n111 DGND.t221 144.886
R488 DGND.n802 DGND.t488 144.886
R489 DGND.n712 DGND.t407 144.886
R490 DGND.n581 DGND.t53 144.886
R491 DGND.n558 DGND.t428 144.886
R492 DGND.n631 DGND.t145 144.886
R493 DGND.n458 DGND.t172 144.886
R494 DGND.n1 DGND.t528 144.886
R495 DGND.n38 DGND.t190 144.886
R496 DGND.n384 DGND.t147 144.886
R497 DGND.n339 DGND.t174 144.886
R498 DGND.n830 DGND.n829 97.1434
R499 DGND.n233 DGND.n232 97.1434
R500 DGND.n515 DGND.n514 97.1434
R501 DGND.n673 DGND.n672 97.1434
R502 DGND.t141 DGND.t474 95.6527
R503 DGND.t203 DGND.t258 95.6527
R504 DGND.t265 DGND.t458 95.6527
R505 DGND.t151 DGND.t321 95.6527
R506 DGND.t497 DGND.t306 88.2948
R507 DGND.t280 DGND.t462 88.2948
R508 DGND.t385 DGND.t175 88.2948
R509 DGND.t512 DGND.t98 88.2948
R510 DGND.t476 DGND.t25 88.2948
R511 DGND.t73 DGND.t112 88.2948
R512 DGND.t19 DGND.t229 88.2948
R513 DGND.t414 DGND.t475 88.2948
R514 DGND.n820 DGND.t155 74.2862
R515 DGND.n88 DGND.t197 74.2862
R516 DGND.n612 DGND.t364 74.2862
R517 DGND.n615 DGND.t455 74.2862
R518 DGND.t317 DGND.t535 66.2212
R519 DGND.t237 DGND.t159 66.2212
R520 DGND.t33 DGND.t194 66.2212
R521 DGND.t200 DGND.t408 66.2212
R522 DGND.t525 DGND.t339 66.2212
R523 DGND.t377 DGND.t319 66.2212
R524 DGND.t350 DGND.t26 66.2212
R525 DGND.t93 DGND.t446 66.2212
R526 DGND.n829 DGND.t5 61.4291
R527 DGND.n233 DGND.t224 61.4291
R528 DGND.n515 DGND.t358 61.4291
R529 DGND.n673 DGND.t507 61.4291
R530 DGND.t370 DGND.t417 44.1477
R531 DGND.t142 DGND.t337 44.1477
R532 DGND.t186 DGND.t372 44.1477
R533 DGND.t465 DGND.t284 44.1477
R534 DGND.t481 DGND.t282 44.1477
R535 DGND.t274 DGND.t450 44.1477
R536 DGND.t184 DGND.t513 44.1477
R537 DGND.t31 DGND.t43 44.1477
R538 DGND.t367 DGND.t387 44.1477
R539 DGND.t368 DGND.t344 44.1477
R540 DGND.t359 DGND.t257 44.1477
R541 DGND.t288 DGND.t499 44.1477
R542 DGND.t97 DGND.t389 44.1477
R543 DGND.t132 DGND.t342 44.1477
R544 DGND.t176 DGND.t431 44.1477
R545 DGND.t6 DGND.t439 44.1477
R546 DGND.t502 DGND.t252 44.1477
R547 DGND.t437 DGND.t384 44.1477
R548 DGND.t480 DGND.t435 44.1477
R549 DGND.t264 DGND.t82 44.1477
R550 DGND.t39 DGND.t537 44.1477
R551 DGND.t419 DGND.t108 44.1477
R552 DGND.t148 DGND.t421 44.1477
R553 DGND.t193 DGND.t425 44.1477
R554 DGND.n77 DGND.n76 43.9358
R555 DGND.n871 DGND.n870 43.9358
R556 DGND.n879 DGND.n878 43.9358
R557 DGND.n244 DGND.n243 43.9358
R558 DGND.n252 DGND.n251 43.9358
R559 DGND.n307 DGND.n305 43.9358
R560 DGND.n148 DGND.n147 43.9358
R561 DGND.n185 DGND.n184 43.9358
R562 DGND.n193 DGND.n192 43.9358
R563 DGND.n775 DGND.n774 43.9358
R564 DGND.n783 DGND.n782 43.9358
R565 DGND.n735 DGND.n702 43.9358
R566 DGND.n597 DGND.n596 43.9358
R567 DGND.n537 DGND.n536 43.9358
R568 DGND.n526 DGND.n525 43.9358
R569 DGND.n669 DGND.n620 43.9358
R570 DGND.n660 DGND.n623 43.9358
R571 DGND.n478 DGND.n476 43.9358
R572 DGND.n962 DGND.n961 43.9358
R573 DGND.n931 DGND.n930 43.9358
R574 DGND.n939 DGND.n938 43.9358
R575 DGND.n429 DGND.n17 43.9358
R576 DGND.n418 DGND.n417 43.9358
R577 DGND.n409 DGND.n408 43.9358
R578 DGND.n359 DGND.n357 43.9358
R579 DGND.n45 DGND.t195 38.5719
R580 DGND.n45 DGND.t210 38.5719
R581 DGND.n50 DGND.t411 38.5719
R582 DGND.n50 DGND.t226 38.5719
R583 DGND.n833 DGND.t89 38.5719
R584 DGND.n833 DGND.t29 38.5719
R585 DGND.n838 DGND.t294 38.5719
R586 DGND.n838 DGND.t185 38.5719
R587 DGND.n216 DGND.t275 38.5719
R588 DGND.n216 DGND.t464 38.5719
R589 DGND.n223 DGND.t484 38.5719
R590 DGND.n223 DGND.t279 38.5719
R591 DGND.n279 DGND.t56 38.5719
R592 DGND.n279 DGND.t81 38.5719
R593 DGND.n275 DGND.t269 38.5719
R594 DGND.n275 DGND.t160 38.5719
R595 DGND.n830 DGND.t153 38.5719
R596 DGND.n232 DGND.t199 38.5719
R597 DGND.n116 DGND.t536 38.5719
R598 DGND.n116 DGND.t219 38.5719
R599 DGND.n121 DGND.t131 38.5719
R600 DGND.n121 DGND.t240 38.5719
R601 DGND.n97 DGND.t479 38.5719
R602 DGND.n97 DGND.t140 38.5719
R603 DGND.n102 DGND.t297 38.5719
R604 DGND.n102 DGND.t371 38.5719
R605 DGND.n751 DGND.t500 38.5719
R606 DGND.n751 DGND.t541 38.5719
R607 DGND.n758 DGND.t260 38.5719
R608 DGND.n758 DGND.t516 38.5719
R609 DGND.n723 DGND.t111 38.5719
R610 DGND.n723 DGND.t22 38.5719
R611 DGND.n730 DGND.t59 38.5719
R612 DGND.n730 DGND.t409 38.5719
R613 DGND.n564 DGND.t320 38.5719
R614 DGND.n564 DGND.t2 38.5719
R615 DGND.n570 DGND.t127 38.5719
R616 DGND.n570 DGND.t392 38.5719
R617 DGND.n530 DGND.t332 38.5719
R618 DGND.n530 DGND.t250 38.5719
R619 DGND.n541 DGND.t509 38.5719
R620 DGND.n541 DGND.t440 38.5719
R621 DGND.n642 DGND.t177 38.5719
R622 DGND.n642 DGND.t120 38.5719
R623 DGND.n655 DGND.t135 38.5719
R624 DGND.n655 DGND.t254 38.5719
R625 DGND.n450 DGND.t348 38.5719
R626 DGND.n450 DGND.t486 38.5719
R627 DGND.n446 DGND.t205 38.5719
R628 DGND.n446 DGND.t340 38.5719
R629 DGND.n514 DGND.t362 38.5719
R630 DGND.n672 DGND.t457 38.5719
R631 DGND.n8 DGND.t447 38.5719
R632 DGND.n8 DGND.t346 38.5719
R633 DGND.n967 DGND.t42 38.5719
R634 DGND.n967 DGND.t494 38.5719
R635 DGND.n24 DGND.t445 38.5719
R636 DGND.n24 DGND.t150 38.5719
R637 DGND.n29 DGND.t413 38.5719
R638 DGND.n29 DGND.t420 38.5719
R639 DGND.n401 DGND.t40 38.5719
R640 DGND.n401 DGND.t520 38.5719
R641 DGND.n374 DGND.t267 38.5719
R642 DGND.n374 DGND.t434 38.5719
R643 DGND.n331 DGND.t313 38.5719
R644 DGND.n331 DGND.t122 38.5719
R645 DGND.n327 DGND.t402 38.5719
R646 DGND.n327 DGND.t27 38.5719
R647 DGND.n897 DGND.n43 34.6358
R648 DGND.n81 DGND.n43 34.6358
R649 DGND.n81 DGND.n80 34.6358
R650 DGND.n72 DGND.n71 34.6358
R651 DGND.n68 DGND.n67 34.6358
R652 DGND.n67 DGND.n66 34.6358
R653 DGND.n66 DGND.n57 34.6358
R654 DGND.n882 DGND.n826 34.6358
R655 DGND.n876 DGND.n826 34.6358
R656 DGND.n876 DGND.n875 34.6358
R657 DGND.n866 DGND.n865 34.6358
R658 DGND.n863 DGND.n839 34.6358
R659 DGND.n855 DGND.n839 34.6358
R660 DGND.n855 DGND.n854 34.6358
R661 DGND.n266 DGND.n265 34.6358
R662 DGND.n265 DGND.n212 34.6358
R663 DGND.n257 DGND.n212 34.6358
R664 DGND.n255 DGND.n217 34.6358
R665 DGND.n247 DGND.n224 34.6358
R666 DGND.n228 DGND.n224 34.6358
R667 DGND.n240 DGND.n228 34.6358
R668 DGND.n291 DGND.n290 34.6358
R669 DGND.n293 DGND.n291 34.6358
R670 DGND.n293 DGND.n292 34.6358
R671 DGND.n301 DGND.n300 34.6358
R672 DGND.n311 DGND.n310 34.6358
R673 DGND.n311 DGND.n273 34.6358
R674 DGND.n319 DGND.n273 34.6358
R675 DGND.n59 DGND.n58 34.6358
R676 DGND.n60 DGND.n59 34.6358
R677 DGND.n851 DGND.n843 34.6358
R678 DGND.n851 DGND.n850 34.6358
R679 DGND.n888 DGND.n822 34.6358
R680 DGND.n888 DGND.n887 34.6358
R681 DGND.n887 DGND.n886 34.6358
R682 DGND.n236 DGND.n235 34.6358
R683 DGND.n236 DGND.n89 34.6358
R684 DGND.n816 DGND.n89 34.6358
R685 DGND.n270 DGND.n269 34.6358
R686 DGND.n269 DGND.n208 34.6358
R687 DGND.n288 DGND.n283 34.6358
R688 DGND.n295 DGND.n283 34.6358
R689 DGND.n159 DGND.n113 34.6358
R690 DGND.n152 DGND.n113 34.6358
R691 DGND.n152 DGND.n151 34.6358
R692 DGND.n143 DGND.n142 34.6358
R693 DGND.n139 DGND.n138 34.6358
R694 DGND.n138 DGND.n137 34.6358
R695 DGND.n137 DGND.n128 34.6358
R696 DGND.n196 DGND.n94 34.6358
R697 DGND.n190 DGND.n94 34.6358
R698 DGND.n190 DGND.n189 34.6358
R699 DGND.n180 DGND.n179 34.6358
R700 DGND.n177 DGND.n103 34.6358
R701 DGND.n169 DGND.n103 34.6358
R702 DGND.n169 DGND.n168 34.6358
R703 DGND.n797 DGND.n796 34.6358
R704 DGND.n796 DGND.n747 34.6358
R705 DGND.n788 DGND.n747 34.6358
R706 DGND.n786 DGND.n752 34.6358
R707 DGND.n778 DGND.n759 34.6358
R708 DGND.n763 DGND.n759 34.6358
R709 DGND.n771 DGND.n763 34.6358
R710 DGND.n716 DGND.n715 34.6358
R711 DGND.n716 DGND.n706 34.6358
R712 DGND.n722 DGND.n706 34.6358
R713 DGND.n726 DGND.n725 34.6358
R714 DGND.n731 DGND.n700 34.6358
R715 DGND.n740 DGND.n700 34.6358
R716 DGND.n741 DGND.n740 34.6358
R717 DGND.n130 DGND.n129 34.6358
R718 DGND.n131 DGND.n130 34.6358
R719 DGND.n165 DGND.n107 34.6358
R720 DGND.n165 DGND.n164 34.6358
R721 DGND.n200 DGND.n92 34.6358
R722 DGND.n193 DGND.n92 34.6358
R723 DGND.n774 DGND.n761 34.6358
R724 DGND.n766 DGND.n761 34.6358
R725 DGND.n801 DGND.n800 34.6358
R726 DGND.n800 DGND.n743 34.6358
R727 DGND.n718 DGND.n710 34.6358
R728 DGND.n719 DGND.n718 34.6358
R729 DGND.n602 DGND.n563 34.6358
R730 DGND.n602 DGND.n601 34.6358
R731 DGND.n601 DGND.n600 34.6358
R732 DGND.n592 DGND.n591 34.6358
R733 DGND.n588 DGND.n587 34.6358
R734 DGND.n587 DGND.n586 34.6358
R735 DGND.n586 DGND.n577 34.6358
R736 DGND.n522 DGND.n521 34.6358
R737 DGND.n521 DGND.n506 34.6358
R738 DGND.n529 DGND.n506 34.6358
R739 DGND.n540 DGND.n502 34.6358
R740 DGND.n543 DGND.n497 34.6358
R741 DGND.n551 DGND.n497 34.6358
R742 DGND.n552 DGND.n551 34.6358
R743 DGND.n641 DGND.n629 34.6358
R744 DGND.n645 DGND.n641 34.6358
R745 DGND.n645 DGND.n644 34.6358
R746 DGND.n653 DGND.n624 34.6358
R747 DGND.n665 DGND.n621 34.6358
R748 DGND.n666 DGND.n665 34.6358
R749 DGND.n666 DGND.n618 34.6358
R750 DGND.n462 DGND.n461 34.6358
R751 DGND.n464 DGND.n462 34.6358
R752 DGND.n464 DGND.n463 34.6358
R753 DGND.n472 DGND.n471 34.6358
R754 DGND.n482 DGND.n481 34.6358
R755 DGND.n482 DGND.n444 34.6358
R756 DGND.n693 DGND.n444 34.6358
R757 DGND.n579 DGND.n578 34.6358
R758 DGND.n580 DGND.n579 34.6358
R759 DGND.n556 DGND.n495 34.6358
R760 DGND.n557 DGND.n556 34.6358
R761 DGND.n611 DGND.n489 34.6358
R762 DGND.n512 DGND.n489 34.6358
R763 DGND.n517 DGND.n512 34.6358
R764 DGND.n671 DGND.n616 34.6358
R765 DGND.n682 DGND.n616 34.6358
R766 DGND.n683 DGND.n682 34.6358
R767 DGND.n637 DGND.n632 34.6358
R768 DGND.n638 DGND.n637 34.6358
R769 DGND.n459 DGND.n454 34.6358
R770 DGND.n466 DGND.n454 34.6358
R771 DGND.n905 DGND.n13 34.6358
R772 DGND.n957 DGND.n13 34.6358
R773 DGND.n958 DGND.n957 34.6358
R774 DGND.n970 DGND.n966 34.6358
R775 DGND.n968 DGND.n2 34.6358
R776 DGND.n978 DGND.n2 34.6358
R777 DGND.n979 DGND.n978 34.6358
R778 DGND.n942 DGND.n21 34.6358
R779 DGND.n936 DGND.n21 34.6358
R780 DGND.n936 DGND.n935 34.6358
R781 DGND.n926 DGND.n925 34.6358
R782 DGND.n923 DGND.n30 34.6358
R783 DGND.n915 DGND.n30 34.6358
R784 DGND.n915 DGND.n914 34.6358
R785 DGND.n391 DGND.n390 34.6358
R786 DGND.n391 DGND.n377 34.6358
R787 DGND.n400 DGND.n377 34.6358
R788 DGND.n405 DGND.n403 34.6358
R789 DGND.n415 DGND.n414 34.6358
R790 DGND.n415 DGND.n370 34.6358
R791 DGND.n421 DGND.n370 34.6358
R792 DGND.n343 DGND.n342 34.6358
R793 DGND.n345 DGND.n343 34.6358
R794 DGND.n345 DGND.n344 34.6358
R795 DGND.n353 DGND.n352 34.6358
R796 DGND.n363 DGND.n362 34.6358
R797 DGND.n363 DGND.n325 34.6358
R798 DGND.n438 DGND.n325 34.6358
R799 DGND.n976 DGND.n974 34.6358
R800 DGND.n976 DGND.n975 34.6358
R801 DGND.n911 DGND.n34 34.6358
R802 DGND.n911 DGND.n910 34.6358
R803 DGND.n946 DGND.n19 34.6358
R804 DGND.n939 DGND.n19 34.6358
R805 DGND.n418 DGND.n368 34.6358
R806 DGND.n425 DGND.n368 34.6358
R807 DGND.n385 DGND.n382 34.6358
R808 DGND.n394 DGND.n382 34.6358
R809 DGND.n340 DGND.n335 34.6358
R810 DGND.n347 DGND.n335 34.6358
R811 DGND.n74 DGND.n46 32.7534
R812 DGND.n874 DGND.n873 32.7534
R813 DGND.n248 DGND.n222 32.7534
R814 DGND.n303 DGND.n276 32.7534
R815 DGND.n145 DGND.n117 32.7534
R816 DGND.n188 DGND.n187 32.7534
R817 DGND.n779 DGND.n757 32.7534
R818 DGND.n732 DGND.n729 32.7534
R819 DGND.n594 DGND.n565 32.7534
R820 DGND.n533 DGND.n532 32.7534
R821 DGND.n657 DGND.n656 32.7534
R822 DGND.n474 DGND.n447 32.7534
R823 DGND.n964 DGND.n9 32.7534
R824 DGND.n934 DGND.n933 32.7534
R825 DGND.n413 DGND.n373 32.7534
R826 DGND.n355 DGND.n328 32.7534
R827 DGND.n898 DGND.n41 29.6299
R828 DGND.n883 DGND.n824 29.6299
R829 DGND.n239 DGND.n238 29.6299
R830 DGND.n321 DGND.n320 29.6299
R831 DGND.n161 DGND.n160 29.6299
R832 DGND.n197 DGND.n91 29.6299
R833 DGND.n770 DGND.n769 29.6299
R834 DGND.n805 DGND.n804 29.6299
R835 DGND.n562 DGND.n560 29.6299
R836 DGND.n520 DGND.n510 29.6299
R837 DGND.n679 DGND.n678 29.6299
R838 DGND.n695 DGND.n694 29.6299
R839 DGND.n907 DGND.n906 29.6299
R840 DGND.n943 DGND.n18 29.6299
R841 DGND.n422 DGND.n367 29.6299
R842 DGND.n440 DGND.n439 29.6299
R843 DGND.n156 DGND.n114 26.6181
R844 DGND.n157 DGND.n156 26.6181
R845 DGND.n891 DGND.n84 26.6181
R846 DGND.n891 DGND.n890 26.6181
R847 DGND.n814 DGND.n813 26.6181
R848 DGND.n813 DGND.n87 26.6181
R849 DGND.n894 DGND.n42 26.6181
R850 DGND.n895 DGND.n894 26.6181
R851 DGND.n316 DGND.n314 26.6181
R852 DGND.n317 DGND.n316 26.6181
R853 DGND.n808 DGND.n204 26.6181
R854 DGND.n808 DGND.n807 26.6181
R855 DGND.n608 DGND.n488 26.6181
R856 DGND.n609 DGND.n608 26.6181
R857 DGND.n687 DGND.n486 26.6181
R858 DGND.n687 DGND.n686 26.6181
R859 DGND.n605 DGND.n491 26.6181
R860 DGND.n605 DGND.n604 26.6181
R861 DGND.n690 DGND.n485 26.6181
R862 DGND.n691 DGND.n690 26.6181
R863 DGND.n950 DGND.n16 26.6181
R864 DGND.n950 DGND.n949 26.6181
R865 DGND.n953 DGND.n15 26.6181
R866 DGND.n954 DGND.n953 26.6181
R867 DGND.n435 DGND.n366 26.6181
R868 DGND.n436 DGND.n435 26.6181
R869 DGND.n820 DGND.t63 25.4291
R870 DGND.n88 DGND.t326 25.4291
R871 DGND.n612 DGND.t125 25.4291
R872 DGND.n615 DGND.t382 25.4291
R873 DGND.n54 DGND.t77 24.9236
R874 DGND.n54 DGND.t165 24.9236
R875 DGND.n858 DGND.t44 24.9236
R876 DGND.n858 DGND.t388 24.9236
R877 DGND.n261 DGND.t285 24.9236
R878 DGND.n261 DGND.t283 24.9236
R879 DGND.n282 DGND.t107 24.9236
R880 DGND.n282 DGND.t67 24.9236
R881 DGND.n125 DGND.t228 24.9236
R882 DGND.n125 DGND.t522 24.9236
R883 DGND.n172 DGND.t338 24.9236
R884 DGND.n172 DGND.t373 24.9236
R885 DGND.n792 DGND.t369 24.9236
R886 DGND.n792 DGND.t360 24.9236
R887 DGND.n709 DGND.t79 24.9236
R888 DGND.n709 DGND.t38 24.9236
R889 DGND.n574 DGND.t394 24.9236
R890 DGND.n574 DGND.t49 24.9236
R891 DGND.n499 DGND.t503 24.9236
R892 DGND.n499 DGND.t438 24.9236
R893 DGND.n626 DGND.t390 24.9236
R894 DGND.n626 DGND.t343 24.9236
R895 DGND.n453 DGND.t492 24.9236
R896 DGND.n453 DGND.t396 24.9236
R897 DGND.n5 DGND.t449 24.9236
R898 DGND.n5 DGND.t46 24.9236
R899 DGND.n918 DGND.t422 24.9236
R900 DGND.n918 DGND.t426 24.9236
R901 DGND.n381 DGND.t436 24.9236
R902 DGND.n381 DGND.t83 24.9236
R903 DGND.n334 DGND.t13 24.9236
R904 DGND.n334 DGND.t300 24.9236
R905 DGND.n898 DGND.n897 24.0946
R906 DGND.n883 DGND.n882 24.0946
R907 DGND.n240 DGND.n239 24.0946
R908 DGND.n320 DGND.n319 24.0946
R909 DGND.n160 DGND.n159 24.0946
R910 DGND.n197 DGND.n196 24.0946
R911 DGND.n771 DGND.n770 24.0946
R912 DGND.n805 DGND.n741 24.0946
R913 DGND.n563 DGND.n562 24.0946
R914 DGND.n522 DGND.n520 24.0946
R915 DGND.n678 DGND.n618 24.0946
R916 DGND.n694 DGND.n693 24.0946
R917 DGND.n906 DGND.n905 24.0946
R918 DGND.n943 DGND.n942 24.0946
R919 DGND.n422 DGND.n421 24.0946
R920 DGND.n439 DGND.n438 24.0946
R921 DGND.n61 DGND.n60 23.7181
R922 DGND.n850 DGND.n847 23.7181
R923 DGND.n271 DGND.n270 23.7181
R924 DGND.n288 DGND.n287 23.7181
R925 DGND.n132 DGND.n131 23.7181
R926 DGND.n164 DGND.n111 23.7181
R927 DGND.n802 DGND.n801 23.7181
R928 DGND.n712 DGND.n710 23.7181
R929 DGND.n581 DGND.n580 23.7181
R930 DGND.n558 DGND.n557 23.7181
R931 DGND.n632 DGND.n631 23.7181
R932 DGND.n459 DGND.n458 23.7181
R933 DGND.n975 DGND.n1 23.7181
R934 DGND.n910 DGND.n38 23.7181
R935 DGND.n385 DGND.n384 23.7181
R936 DGND.n340 DGND.n339 23.7181
R937 DGND.n58 DGND.n55 22.9652
R938 DGND.n859 DGND.n843 22.9652
R939 DGND.n822 DGND.n821 22.9652
R940 DGND.n817 DGND.n816 22.9652
R941 DGND.n262 DGND.n208 22.9652
R942 DGND.n296 DGND.n295 22.9652
R943 DGND.n129 DGND.n126 22.9652
R944 DGND.n173 DGND.n107 22.9652
R945 DGND.n793 DGND.n743 22.9652
R946 DGND.n720 DGND.n719 22.9652
R947 DGND.n578 DGND.n575 22.9652
R948 DGND.n547 DGND.n495 22.9652
R949 DGND.n613 DGND.n611 22.9652
R950 DGND.n684 DGND.n683 22.9652
R951 DGND.n638 DGND.n627 22.9652
R952 DGND.n467 DGND.n466 22.9652
R953 DGND.n974 DGND.n973 22.9652
R954 DGND.n919 DGND.n34 22.9652
R955 DGND.n395 DGND.n394 22.9652
R956 DGND.n348 DGND.n347 22.9652
R957 DGND.n886 DGND.n823 22.2496
R958 DGND.n235 DGND.n234 22.2496
R959 DGND.n517 DGND.n516 22.2496
R960 DGND.n674 DGND.n671 22.2496
R961 DGND.n55 DGND.n53 21.4593
R962 DGND.n860 DGND.n859 21.4593
R963 DGND.n262 DGND.n260 21.4593
R964 DGND.n298 DGND.n296 21.4593
R965 DGND.n126 DGND.n124 21.4593
R966 DGND.n174 DGND.n173 21.4593
R967 DGND.n793 DGND.n791 21.4593
R968 DGND.n720 DGND.n708 21.4593
R969 DGND.n575 DGND.n573 21.4593
R970 DGND.n547 DGND.n546 21.4593
R971 DGND.n648 DGND.n627 21.4593
R972 DGND.n469 DGND.n467 21.4593
R973 DGND.n973 DGND.n972 21.4593
R974 DGND.n920 DGND.n919 21.4593
R975 DGND.n396 DGND.n395 21.4593
R976 DGND.n350 DGND.n348 21.4593
R977 DGND.n201 DGND.n200 19.9534
R978 DGND.n767 DGND.n766 19.9534
R979 DGND.n947 DGND.n946 19.9534
R980 DGND.n426 DGND.n425 19.9534
R981 DGND.n53 DGND.n52 16.9417
R982 DGND.n860 DGND.n842 16.9417
R983 DGND.n260 DGND.n214 16.9417
R984 DGND.n298 DGND.n297 16.9417
R985 DGND.n124 DGND.n123 16.9417
R986 DGND.n174 DGND.n106 16.9417
R987 DGND.n791 DGND.n749 16.9417
R988 DGND.n708 DGND.n705 16.9417
R989 DGND.n573 DGND.n572 16.9417
R990 DGND.n546 DGND.n500 16.9417
R991 DGND.n649 DGND.n648 16.9417
R992 DGND.n469 DGND.n468 16.9417
R993 DGND.n972 DGND.n6 16.9417
R994 DGND.n920 DGND.n33 16.9417
R995 DGND.n397 DGND.n396 16.9417
R996 DGND.n350 DGND.n349 16.9417
R997 DGND.n63 DGND.n62 16.077
R998 DGND.n846 DGND.n845 16.077
R999 DGND.n211 DGND.n209 16.077
R1000 DGND.n286 DGND.n285 16.077
R1001 DGND.n48 DGND.n44 16.077
R1002 DGND.n869 DGND.n868 16.077
R1003 DGND.n220 DGND.n219 16.077
R1004 DGND.n306 DGND.n274 16.077
R1005 DGND.n134 DGND.n133 16.077
R1006 DGND.n110 DGND.n109 16.077
R1007 DGND.n746 DGND.n744 16.077
R1008 DGND.n714 DGND.n713 16.077
R1009 DGND.n119 DGND.n115 16.077
R1010 DGND.n183 DGND.n182 16.077
R1011 DGND.n755 DGND.n754 16.077
R1012 DGND.n737 DGND.n736 16.077
R1013 DGND.n583 DGND.n582 16.077
R1014 DGND.n554 DGND.n553 16.077
R1015 DGND.n635 DGND.n634 16.077
R1016 DGND.n457 DGND.n456 16.077
R1017 DGND.n568 DGND.n566 16.077
R1018 DGND.n505 DGND.n504 16.077
R1019 DGND.n662 DGND.n661 16.077
R1020 DGND.n477 DGND.n445 16.077
R1021 DGND.n981 DGND.n980 16.077
R1022 DGND.n37 DGND.n36 16.077
R1023 DGND.n389 DGND.n388 16.077
R1024 DGND.n338 DGND.n337 16.077
R1025 DGND.n12 DGND.n11 16.077
R1026 DGND.n929 DGND.n928 16.077
R1027 DGND.n431 DGND.n430 16.077
R1028 DGND.n411 DGND.n410 16.077
R1029 DGND.n358 DGND.n326 16.077
R1030 DGND.n879 DGND.n831 11.7085
R1031 DGND.n243 DGND.n226 11.7085
R1032 DGND.n525 DGND.n508 11.7085
R1033 DGND.n670 DGND.n669 11.7085
R1034 DGND.n80 DGND.n46 11.6711
R1035 DGND.n875 DGND.n874 11.6711
R1036 DGND.n248 DGND.n247 11.6711
R1037 DGND.n310 DGND.n276 11.6711
R1038 DGND.n151 DGND.n117 11.6711
R1039 DGND.n189 DGND.n188 11.6711
R1040 DGND.n779 DGND.n778 11.6711
R1041 DGND.n732 DGND.n731 11.6711
R1042 DGND.n600 DGND.n565 11.6711
R1043 DGND.n533 DGND.n529 11.6711
R1044 DGND.n656 DGND.n621 11.6711
R1045 DGND.n481 DGND.n447 11.6711
R1046 DGND.n958 DGND.n9 11.6711
R1047 DGND.n935 DGND.n934 11.6711
R1048 DGND.n414 DGND.n413 11.6711
R1049 DGND.n362 DGND.n328 11.6711
R1050 DGND.n77 DGND.n48 10.5417
R1051 DGND.n870 DGND.n869 10.5417
R1052 DGND.n251 DGND.n219 10.5417
R1053 DGND.n307 DGND.n306 10.5417
R1054 DGND.n148 DGND.n119 10.5417
R1055 DGND.n184 DGND.n183 10.5417
R1056 DGND.n782 DGND.n754 10.5417
R1057 DGND.n736 DGND.n735 10.5417
R1058 DGND.n597 DGND.n568 10.5417
R1059 DGND.n536 DGND.n504 10.5417
R1060 DGND.n661 DGND.n660 10.5417
R1061 DGND.n478 DGND.n477 10.5417
R1062 DGND.n961 DGND.n11 10.5417
R1063 DGND.n930 DGND.n929 10.5417
R1064 DGND.n430 DGND.n429 10.5417
R1065 DGND.n410 DGND.n409 10.5417
R1066 DGND.n359 DGND.n358 10.5417
R1067 DGND.n713 DGND.n712 9.3005
R1068 DGND.n711 DGND.n710 9.3005
R1069 DGND.n718 DGND.n717 9.3005
R1070 DGND.n719 DGND.n707 9.3005
R1071 DGND.n721 DGND.n720 9.3005
R1072 DGND.n708 DGND.n704 9.3005
R1073 DGND.n727 DGND.n705 9.3005
R1074 DGND.n735 DGND.n734 9.3005
R1075 DGND.n803 DGND.n802 9.3005
R1076 DGND.n801 DGND.n742 9.3005
R1077 DGND.n800 DGND.n799 9.3005
R1078 DGND.n745 DGND.n743 9.3005
R1079 DGND.n794 DGND.n793 9.3005
R1080 DGND.n791 DGND.n790 9.3005
R1081 DGND.n750 DGND.n749 9.3005
R1082 DGND.n782 DGND.n781 9.3005
R1083 DGND.n774 DGND.n773 9.3005
R1084 DGND.n762 DGND.n761 9.3005
R1085 DGND.n766 DGND.n765 9.3005
R1086 DGND.n768 DGND.n767 9.3005
R1087 DGND.n202 DGND.n201 9.3005
R1088 DGND.n200 DGND.n199 9.3005
R1089 DGND.n93 DGND.n92 9.3005
R1090 DGND.n194 DGND.n193 9.3005
R1091 DGND.n184 DGND.n100 9.3005
R1092 DGND.n106 DGND.n104 9.3005
R1093 DGND.n175 DGND.n174 9.3005
R1094 DGND.n173 DGND.n171 9.3005
R1095 DGND.n108 DGND.n107 9.3005
R1096 DGND.n166 DGND.n165 9.3005
R1097 DGND.n164 DGND.n163 9.3005
R1098 DGND.n162 DGND.n111 9.3005
R1099 DGND.n149 DGND.n148 9.3005
R1100 DGND.n123 DGND.n120 9.3005
R1101 DGND.n141 DGND.n124 9.3005
R1102 DGND.n140 DGND.n126 9.3005
R1103 DGND.n129 DGND.n127 9.3005
R1104 DGND.n136 DGND.n130 9.3005
R1105 DGND.n135 DGND.n131 9.3005
R1106 DGND.n134 DGND.n132 9.3005
R1107 DGND.n806 DGND.n805 9.3005
R1108 DGND.n715 DGND.n711 9.3005
R1109 DGND.n717 DGND.n716 9.3005
R1110 DGND.n707 DGND.n706 9.3005
R1111 DGND.n722 DGND.n721 9.3005
R1112 DGND.n725 DGND.n704 9.3005
R1113 DGND.n727 DGND.n726 9.3005
R1114 DGND.n729 DGND.n728 9.3005
R1115 DGND.n733 DGND.n732 9.3005
R1116 DGND.n731 DGND.n701 9.3005
R1117 DGND.n738 DGND.n700 9.3005
R1118 DGND.n740 DGND.n739 9.3005
R1119 DGND.n741 DGND.n205 9.3005
R1120 DGND.n770 DGND.n764 9.3005
R1121 DGND.n798 DGND.n797 9.3005
R1122 DGND.n796 DGND.n795 9.3005
R1123 DGND.n748 DGND.n747 9.3005
R1124 DGND.n789 DGND.n788 9.3005
R1125 DGND.n786 DGND.n785 9.3005
R1126 DGND.n784 DGND.n752 9.3005
R1127 DGND.n757 DGND.n753 9.3005
R1128 DGND.n780 DGND.n779 9.3005
R1129 DGND.n778 DGND.n777 9.3005
R1130 DGND.n776 DGND.n759 9.3005
R1131 DGND.n763 DGND.n760 9.3005
R1132 DGND.n772 DGND.n771 9.3005
R1133 DGND.n198 DGND.n197 9.3005
R1134 DGND.n196 DGND.n195 9.3005
R1135 DGND.n95 DGND.n94 9.3005
R1136 DGND.n191 DGND.n190 9.3005
R1137 DGND.n189 DGND.n96 9.3005
R1138 DGND.n188 DGND.n98 9.3005
R1139 DGND.n187 DGND.n186 9.3005
R1140 DGND.n181 DGND.n180 9.3005
R1141 DGND.n179 DGND.n101 9.3005
R1142 DGND.n177 DGND.n176 9.3005
R1143 DGND.n105 DGND.n103 9.3005
R1144 DGND.n170 DGND.n169 9.3005
R1145 DGND.n168 DGND.n167 9.3005
R1146 DGND.n160 DGND.n112 9.3005
R1147 DGND.n159 DGND.n158 9.3005
R1148 DGND.n154 DGND.n113 9.3005
R1149 DGND.n153 DGND.n152 9.3005
R1150 DGND.n151 DGND.n150 9.3005
R1151 DGND.n118 DGND.n117 9.3005
R1152 DGND.n146 DGND.n145 9.3005
R1153 DGND.n143 DGND.n120 9.3005
R1154 DGND.n142 DGND.n141 9.3005
R1155 DGND.n140 DGND.n139 9.3005
R1156 DGND.n138 DGND.n127 9.3005
R1157 DGND.n137 DGND.n136 9.3005
R1158 DGND.n135 DGND.n128 9.3005
R1159 DGND.n458 DGND.n457 9.3005
R1160 DGND.n460 DGND.n459 9.3005
R1161 DGND.n455 DGND.n454 9.3005
R1162 DGND.n466 DGND.n465 9.3005
R1163 DGND.n467 DGND.n452 9.3005
R1164 DGND.n470 DGND.n469 9.3005
R1165 DGND.n468 DGND.n449 9.3005
R1166 DGND.n479 DGND.n478 9.3005
R1167 DGND.n631 DGND.n443 9.3005
R1168 DGND.n633 DGND.n632 9.3005
R1169 DGND.n637 DGND.n636 9.3005
R1170 DGND.n639 DGND.n638 9.3005
R1171 DGND.n628 DGND.n627 9.3005
R1172 DGND.n648 DGND.n647 9.3005
R1173 DGND.n650 DGND.n649 9.3005
R1174 DGND.n660 DGND.n659 9.3005
R1175 DGND.n669 DGND.n668 9.3005
R1176 DGND.n676 DGND.n675 9.3005
R1177 DGND.n671 DGND.n617 9.3005
R1178 DGND.n680 DGND.n616 9.3005
R1179 DGND.n682 DGND.n681 9.3005
R1180 DGND.n683 DGND.n487 9.3005
R1181 DGND.n611 DGND.n610 9.3005
R1182 DGND.n490 DGND.n489 9.3005
R1183 DGND.n512 DGND.n511 9.3005
R1184 DGND.n518 DGND.n517 9.3005
R1185 DGND.n513 DGND.n509 9.3005
R1186 DGND.n525 DGND.n524 9.3005
R1187 DGND.n536 DGND.n535 9.3005
R1188 DGND.n501 DGND.n500 9.3005
R1189 DGND.n546 DGND.n545 9.3005
R1190 DGND.n548 DGND.n547 9.3005
R1191 DGND.n549 DGND.n495 9.3005
R1192 DGND.n556 DGND.n555 9.3005
R1193 DGND.n557 DGND.n494 9.3005
R1194 DGND.n559 DGND.n558 9.3005
R1195 DGND.n598 DGND.n597 9.3005
R1196 DGND.n572 DGND.n569 9.3005
R1197 DGND.n590 DGND.n573 9.3005
R1198 DGND.n589 DGND.n575 9.3005
R1199 DGND.n578 DGND.n576 9.3005
R1200 DGND.n585 DGND.n579 9.3005
R1201 DGND.n584 DGND.n580 9.3005
R1202 DGND.n583 DGND.n581 9.3005
R1203 DGND.n694 DGND.n442 9.3005
R1204 DGND.n461 DGND.n460 9.3005
R1205 DGND.n462 DGND.n455 9.3005
R1206 DGND.n465 DGND.n464 9.3005
R1207 DGND.n463 DGND.n452 9.3005
R1208 DGND.n471 DGND.n470 9.3005
R1209 DGND.n472 DGND.n449 9.3005
R1210 DGND.n475 DGND.n474 9.3005
R1211 DGND.n448 DGND.n447 9.3005
R1212 DGND.n481 DGND.n480 9.3005
R1213 DGND.n483 DGND.n482 9.3005
R1214 DGND.n484 DGND.n444 9.3005
R1215 DGND.n693 DGND.n692 9.3005
R1216 DGND.n678 DGND.n677 9.3005
R1217 DGND.n630 DGND.n629 9.3005
R1218 DGND.n641 DGND.n640 9.3005
R1219 DGND.n646 DGND.n645 9.3005
R1220 DGND.n644 DGND.n625 9.3005
R1221 DGND.n651 DGND.n624 9.3005
R1222 DGND.n653 DGND.n652 9.3005
R1223 DGND.n658 DGND.n657 9.3005
R1224 DGND.n656 DGND.n622 9.3005
R1225 DGND.n663 DGND.n621 9.3005
R1226 DGND.n665 DGND.n664 9.3005
R1227 DGND.n667 DGND.n666 9.3005
R1228 DGND.n619 DGND.n618 9.3005
R1229 DGND.n520 DGND.n519 9.3005
R1230 DGND.n523 DGND.n522 9.3005
R1231 DGND.n521 DGND.n507 9.3005
R1232 DGND.n527 DGND.n506 9.3005
R1233 DGND.n529 DGND.n528 9.3005
R1234 DGND.n534 DGND.n533 9.3005
R1235 DGND.n532 DGND.n503 9.3005
R1236 DGND.n538 DGND.n502 9.3005
R1237 DGND.n540 DGND.n539 9.3005
R1238 DGND.n544 DGND.n543 9.3005
R1239 DGND.n498 DGND.n497 9.3005
R1240 DGND.n551 DGND.n550 9.3005
R1241 DGND.n552 DGND.n496 9.3005
R1242 DGND.n562 DGND.n561 9.3005
R1243 DGND.n563 DGND.n492 9.3005
R1244 DGND.n603 DGND.n602 9.3005
R1245 DGND.n601 DGND.n493 9.3005
R1246 DGND.n600 DGND.n599 9.3005
R1247 DGND.n567 DGND.n565 9.3005
R1248 DGND.n595 DGND.n594 9.3005
R1249 DGND.n592 DGND.n569 9.3005
R1250 DGND.n591 DGND.n590 9.3005
R1251 DGND.n589 DGND.n588 9.3005
R1252 DGND.n587 DGND.n576 9.3005
R1253 DGND.n586 DGND.n585 9.3005
R1254 DGND.n584 DGND.n577 9.3005
R1255 DGND.n287 DGND.n286 9.3005
R1256 DGND.n289 DGND.n288 9.3005
R1257 DGND.n284 DGND.n283 9.3005
R1258 DGND.n295 DGND.n294 9.3005
R1259 DGND.n296 DGND.n281 9.3005
R1260 DGND.n299 DGND.n298 9.3005
R1261 DGND.n297 DGND.n278 9.3005
R1262 DGND.n308 DGND.n307 9.3005
R1263 DGND.n272 DGND.n271 9.3005
R1264 DGND.n270 DGND.n207 9.3005
R1265 DGND.n269 DGND.n268 9.3005
R1266 DGND.n210 DGND.n208 9.3005
R1267 DGND.n263 DGND.n262 9.3005
R1268 DGND.n260 DGND.n259 9.3005
R1269 DGND.n215 DGND.n214 9.3005
R1270 DGND.n251 DGND.n250 9.3005
R1271 DGND.n243 DGND.n242 9.3005
R1272 DGND.n231 DGND.n227 9.3005
R1273 DGND.n235 DGND.n230 9.3005
R1274 DGND.n237 DGND.n236 9.3005
R1275 DGND.n90 DGND.n89 9.3005
R1276 DGND.n816 DGND.n815 9.3005
R1277 DGND.n822 DGND.n85 9.3005
R1278 DGND.n889 DGND.n888 9.3005
R1279 DGND.n887 DGND.n86 9.3005
R1280 DGND.n886 DGND.n885 9.3005
R1281 DGND.n828 DGND.n825 9.3005
R1282 DGND.n880 DGND.n879 9.3005
R1283 DGND.n870 DGND.n836 9.3005
R1284 DGND.n842 DGND.n840 9.3005
R1285 DGND.n861 DGND.n860 9.3005
R1286 DGND.n859 DGND.n857 9.3005
R1287 DGND.n844 DGND.n843 9.3005
R1288 DGND.n852 DGND.n851 9.3005
R1289 DGND.n850 DGND.n849 9.3005
R1290 DGND.n848 DGND.n847 9.3005
R1291 DGND.n78 DGND.n77 9.3005
R1292 DGND.n52 DGND.n49 9.3005
R1293 DGND.n70 DGND.n53 9.3005
R1294 DGND.n69 DGND.n55 9.3005
R1295 DGND.n58 DGND.n56 9.3005
R1296 DGND.n65 DGND.n59 9.3005
R1297 DGND.n64 DGND.n60 9.3005
R1298 DGND.n63 DGND.n61 9.3005
R1299 DGND.n320 DGND.n206 9.3005
R1300 DGND.n290 DGND.n289 9.3005
R1301 DGND.n291 DGND.n284 9.3005
R1302 DGND.n294 DGND.n293 9.3005
R1303 DGND.n292 DGND.n281 9.3005
R1304 DGND.n300 DGND.n299 9.3005
R1305 DGND.n301 DGND.n278 9.3005
R1306 DGND.n304 DGND.n303 9.3005
R1307 DGND.n277 DGND.n276 9.3005
R1308 DGND.n310 DGND.n309 9.3005
R1309 DGND.n312 DGND.n311 9.3005
R1310 DGND.n313 DGND.n273 9.3005
R1311 DGND.n319 DGND.n318 9.3005
R1312 DGND.n239 DGND.n229 9.3005
R1313 DGND.n267 DGND.n266 9.3005
R1314 DGND.n265 DGND.n264 9.3005
R1315 DGND.n213 DGND.n212 9.3005
R1316 DGND.n258 DGND.n257 9.3005
R1317 DGND.n255 DGND.n254 9.3005
R1318 DGND.n253 DGND.n217 9.3005
R1319 DGND.n222 DGND.n218 9.3005
R1320 DGND.n249 DGND.n248 9.3005
R1321 DGND.n247 DGND.n246 9.3005
R1322 DGND.n245 DGND.n224 9.3005
R1323 DGND.n228 DGND.n225 9.3005
R1324 DGND.n241 DGND.n240 9.3005
R1325 DGND.n884 DGND.n883 9.3005
R1326 DGND.n882 DGND.n881 9.3005
R1327 DGND.n827 DGND.n826 9.3005
R1328 DGND.n877 DGND.n876 9.3005
R1329 DGND.n875 DGND.n832 9.3005
R1330 DGND.n874 DGND.n834 9.3005
R1331 DGND.n873 DGND.n872 9.3005
R1332 DGND.n867 DGND.n866 9.3005
R1333 DGND.n865 DGND.n837 9.3005
R1334 DGND.n863 DGND.n862 9.3005
R1335 DGND.n841 DGND.n839 9.3005
R1336 DGND.n856 DGND.n855 9.3005
R1337 DGND.n854 DGND.n853 9.3005
R1338 DGND.n899 DGND.n898 9.3005
R1339 DGND.n897 DGND.n896 9.3005
R1340 DGND.n83 DGND.n43 9.3005
R1341 DGND.n82 DGND.n81 9.3005
R1342 DGND.n80 DGND.n79 9.3005
R1343 DGND.n47 DGND.n46 9.3005
R1344 DGND.n75 DGND.n74 9.3005
R1345 DGND.n72 DGND.n49 9.3005
R1346 DGND.n71 DGND.n70 9.3005
R1347 DGND.n69 DGND.n68 9.3005
R1348 DGND.n67 DGND.n56 9.3005
R1349 DGND.n66 DGND.n65 9.3005
R1350 DGND.n64 DGND.n57 9.3005
R1351 DGND.n339 DGND.n338 9.3005
R1352 DGND.n341 DGND.n340 9.3005
R1353 DGND.n336 DGND.n335 9.3005
R1354 DGND.n347 DGND.n346 9.3005
R1355 DGND.n348 DGND.n333 9.3005
R1356 DGND.n351 DGND.n350 9.3005
R1357 DGND.n349 DGND.n330 9.3005
R1358 DGND.n360 DGND.n359 9.3005
R1359 DGND.n384 DGND.n324 9.3005
R1360 DGND.n386 DGND.n385 9.3005
R1361 DGND.n387 DGND.n382 9.3005
R1362 DGND.n394 DGND.n393 9.3005
R1363 DGND.n395 DGND.n380 9.3005
R1364 DGND.n396 DGND.n378 9.3005
R1365 DGND.n398 DGND.n397 9.3005
R1366 DGND.n409 DGND.n375 9.3005
R1367 DGND.n419 DGND.n418 9.3005
R1368 DGND.n369 DGND.n368 9.3005
R1369 DGND.n425 DGND.n424 9.3005
R1370 DGND.n427 DGND.n426 9.3005
R1371 DGND.n429 DGND.n428 9.3005
R1372 DGND.n948 DGND.n947 9.3005
R1373 DGND.n946 DGND.n945 9.3005
R1374 DGND.n20 DGND.n19 9.3005
R1375 DGND.n940 DGND.n939 9.3005
R1376 DGND.n930 DGND.n27 9.3005
R1377 DGND.n33 DGND.n31 9.3005
R1378 DGND.n921 DGND.n920 9.3005
R1379 DGND.n919 DGND.n917 9.3005
R1380 DGND.n35 DGND.n34 9.3005
R1381 DGND.n912 DGND.n911 9.3005
R1382 DGND.n910 DGND.n909 9.3005
R1383 DGND.n908 DGND.n38 9.3005
R1384 DGND.n961 DGND.n960 9.3005
R1385 DGND.n7 DGND.n6 9.3005
R1386 DGND.n972 DGND.n971 9.3005
R1387 DGND.n973 DGND.n4 9.3005
R1388 DGND.n974 DGND.n3 9.3005
R1389 DGND.n977 DGND.n976 9.3005
R1390 DGND.n975 DGND.n0 9.3005
R1391 DGND.n981 DGND.n1 9.3005
R1392 DGND.n439 DGND.n323 9.3005
R1393 DGND.n342 DGND.n341 9.3005
R1394 DGND.n343 DGND.n336 9.3005
R1395 DGND.n346 DGND.n345 9.3005
R1396 DGND.n344 DGND.n333 9.3005
R1397 DGND.n352 DGND.n351 9.3005
R1398 DGND.n353 DGND.n330 9.3005
R1399 DGND.n356 DGND.n355 9.3005
R1400 DGND.n329 DGND.n328 9.3005
R1401 DGND.n362 DGND.n361 9.3005
R1402 DGND.n364 DGND.n363 9.3005
R1403 DGND.n365 DGND.n325 9.3005
R1404 DGND.n438 DGND.n437 9.3005
R1405 DGND.n423 DGND.n422 9.3005
R1406 DGND.n390 DGND.n383 9.3005
R1407 DGND.n392 DGND.n391 9.3005
R1408 DGND.n379 DGND.n377 9.3005
R1409 DGND.n400 DGND.n399 9.3005
R1410 DGND.n403 DGND.n376 9.3005
R1411 DGND.n406 DGND.n405 9.3005
R1412 DGND.n407 DGND.n373 9.3005
R1413 DGND.n413 DGND.n412 9.3005
R1414 DGND.n414 DGND.n372 9.3005
R1415 DGND.n416 DGND.n415 9.3005
R1416 DGND.n371 DGND.n370 9.3005
R1417 DGND.n421 DGND.n420 9.3005
R1418 DGND.n944 DGND.n943 9.3005
R1419 DGND.n942 DGND.n941 9.3005
R1420 DGND.n22 DGND.n21 9.3005
R1421 DGND.n937 DGND.n936 9.3005
R1422 DGND.n935 DGND.n23 9.3005
R1423 DGND.n934 DGND.n25 9.3005
R1424 DGND.n933 DGND.n932 9.3005
R1425 DGND.n927 DGND.n926 9.3005
R1426 DGND.n925 DGND.n28 9.3005
R1427 DGND.n923 DGND.n922 9.3005
R1428 DGND.n32 DGND.n30 9.3005
R1429 DGND.n916 DGND.n915 9.3005
R1430 DGND.n914 DGND.n913 9.3005
R1431 DGND.n906 DGND.n904 9.3005
R1432 DGND.n905 DGND.n14 9.3005
R1433 DGND.n955 DGND.n13 9.3005
R1434 DGND.n957 DGND.n956 9.3005
R1435 DGND.n959 DGND.n958 9.3005
R1436 DGND.n10 DGND.n9 9.3005
R1437 DGND.n964 DGND.n963 9.3005
R1438 DGND.n966 DGND.n7 9.3005
R1439 DGND.n971 DGND.n970 9.3005
R1440 DGND.n968 DGND.n4 9.3005
R1441 DGND.n3 DGND.n2 9.3005
R1442 DGND.n978 DGND.n977 9.3005
R1443 DGND.n979 DGND.n0 9.3005
R1444 DGND.n698 DGND.n322 8.75713
R1445 DGND.n697 DGND.n441 8.75713
R1446 DGND.n903 DGND.n902 8.75713
R1447 DGND.n901 DGND.n900 8.7565
R1448 DGND.n901 DGND.n40 7.91114
R1449 DGND.n902 DGND.n39 7.9105
R1450 DGND.n699 DGND.n698 7.9105
R1451 DGND.n697 DGND.n696 7.9105
R1452 DGND.n71 DGND.n51 7.15344
R1453 DGND.n865 DGND.n864 7.15344
R1454 DGND.n256 DGND.n255 7.15344
R1455 DGND.n300 DGND.n280 7.15344
R1456 DGND.n142 DGND.n122 7.15344
R1457 DGND.n179 DGND.n178 7.15344
R1458 DGND.n787 DGND.n786 7.15344
R1459 DGND.n725 DGND.n724 7.15344
R1460 DGND.n591 DGND.n571 7.15344
R1461 DGND.n542 DGND.n540 7.15344
R1462 DGND.n643 DGND.n624 7.15344
R1463 DGND.n471 DGND.n451 7.15344
R1464 DGND.n970 DGND.n969 7.15344
R1465 DGND.n925 DGND.n924 7.15344
R1466 DGND.n403 DGND.n402 7.15344
R1467 DGND.n352 DGND.n332 7.15344
R1468 DGND.n818 DGND.n817 7.13003
R1469 DGND.n685 DGND.n684 7.13003
R1470 DGND.n614 DGND.n613 7.13003
R1471 DGND.n821 DGND.n819 7.13003
R1472 DGND.n74 DGND.n73 5.64756
R1473 DGND.n873 DGND.n835 5.64756
R1474 DGND.n222 DGND.n221 5.64756
R1475 DGND.n303 DGND.n302 5.64756
R1476 DGND.n145 DGND.n144 5.64756
R1477 DGND.n187 DGND.n99 5.64756
R1478 DGND.n757 DGND.n756 5.64756
R1479 DGND.n729 DGND.n703 5.64756
R1480 DGND.n594 DGND.n593 5.64756
R1481 DGND.n532 DGND.n531 5.64756
R1482 DGND.n657 DGND.n654 5.64756
R1483 DGND.n474 DGND.n473 5.64756
R1484 DGND.n965 DGND.n964 5.64756
R1485 DGND.n933 DGND.n26 5.64756
R1486 DGND.n404 DGND.n373 5.64756
R1487 DGND.n355 DGND.n354 5.64756
R1488 DGND.n831 DGND.n828 4.35795
R1489 DGND.n231 DGND.n226 4.35795
R1490 DGND.n513 DGND.n508 4.35795
R1491 DGND.n675 DGND.n670 4.35795
R1492 DGND.n73 DGND.n72 4.14168
R1493 DGND.n866 DGND.n835 4.14168
R1494 DGND.n221 DGND.n217 4.14168
R1495 DGND.n302 DGND.n301 4.14168
R1496 DGND.n144 DGND.n143 4.14168
R1497 DGND.n180 DGND.n99 4.14168
R1498 DGND.n756 DGND.n752 4.14168
R1499 DGND.n726 DGND.n703 4.14168
R1500 DGND.n593 DGND.n592 4.14168
R1501 DGND.n531 DGND.n502 4.14168
R1502 DGND.n654 DGND.n653 4.14168
R1503 DGND.n473 DGND.n472 4.14168
R1504 DGND.n966 DGND.n965 4.14168
R1505 DGND.n926 DGND.n26 4.14168
R1506 DGND.n405 DGND.n404 4.14168
R1507 DGND.n354 DGND.n353 4.14168
R1508 DGND.n62 DGND.n57 3.01226
R1509 DGND.n854 DGND.n845 3.01226
R1510 DGND.n266 DGND.n211 3.01226
R1511 DGND.n290 DGND.n285 3.01226
R1512 DGND.n133 DGND.n128 3.01226
R1513 DGND.n168 DGND.n109 3.01226
R1514 DGND.n797 DGND.n746 3.01226
R1515 DGND.n715 DGND.n714 3.01226
R1516 DGND.n582 DGND.n577 3.01226
R1517 DGND.n553 DGND.n552 3.01226
R1518 DGND.n634 DGND.n629 3.01226
R1519 DGND.n461 DGND.n456 3.01226
R1520 DGND.n980 DGND.n979 3.01226
R1521 DGND.n914 DGND.n36 3.01226
R1522 DGND.n390 DGND.n389 3.01226
R1523 DGND.n342 DGND.n337 3.01226
R1524 DGND.n68 DGND.n51 2.63579
R1525 DGND.n864 DGND.n863 2.63579
R1526 DGND.n257 DGND.n256 2.63579
R1527 DGND.n292 DGND.n280 2.63579
R1528 DGND.n139 DGND.n122 2.63579
R1529 DGND.n178 DGND.n177 2.63579
R1530 DGND.n788 DGND.n787 2.63579
R1531 DGND.n724 DGND.n722 2.63579
R1532 DGND.n588 DGND.n571 2.63579
R1533 DGND.n543 DGND.n542 2.63579
R1534 DGND.n644 DGND.n643 2.63579
R1535 DGND.n463 DGND.n451 2.63579
R1536 DGND.n969 DGND.n968 2.63579
R1537 DGND.n924 DGND.n923 2.63579
R1538 DGND.n402 DGND.n400 2.63579
R1539 DGND.n344 DGND.n332 2.63579
R1540 DGND.n698 DGND.n697 1.95677
R1541 DGND.n902 DGND.n901 1.86791
R1542 DGND.n828 DGND.n823 1.8161
R1543 DGND.n234 DGND.n231 1.8161
R1544 DGND.n516 DGND.n513 1.8161
R1545 DGND.n675 DGND.n674 1.8161
R1546 DGND.n203 DGND.n202 0.330374
R1547 DGND.n768 DGND.n203 0.330374
R1548 DGND.n432 DGND.n431 0.266946
R1549 DGND.n685 DGND.n614 0.226098
R1550 DGND.n819 DGND.n818 0.226098
R1551 DGND.n432 DGND.n427 0.136132
R1552 DGND.n949 DGND.n948 0.102244
R1553 DGND.n713 DGND.n711 0.0673605
R1554 DGND.n717 DGND.n711 0.0673605
R1555 DGND.n717 DGND.n707 0.0673605
R1556 DGND.n721 DGND.n707 0.0673605
R1557 DGND.n721 DGND.n704 0.0673605
R1558 DGND.n727 DGND.n704 0.0673605
R1559 DGND.n728 DGND.n727 0.0673605
R1560 DGND.n739 DGND.n738 0.0673605
R1561 DGND.n803 DGND.n742 0.0673605
R1562 DGND.n785 DGND.n784 0.0673605
R1563 DGND.n777 DGND.n776 0.0673605
R1564 DGND.n191 DGND.n96 0.0673605
R1565 DGND.n181 DGND.n101 0.0673605
R1566 DGND.n163 DGND.n162 0.0673605
R1567 DGND.n154 DGND.n153 0.0673605
R1568 DGND.n146 DGND.n120 0.0673605
R1569 DGND.n141 DGND.n120 0.0673605
R1570 DGND.n141 DGND.n140 0.0673605
R1571 DGND.n140 DGND.n127 0.0673605
R1572 DGND.n136 DGND.n127 0.0673605
R1573 DGND.n136 DGND.n135 0.0673605
R1574 DGND.n135 DGND.n134 0.0673605
R1575 DGND.n460 DGND.n457 0.0673605
R1576 DGND.n460 DGND.n455 0.0673605
R1577 DGND.n465 DGND.n455 0.0673605
R1578 DGND.n465 DGND.n452 0.0673605
R1579 DGND.n470 DGND.n452 0.0673605
R1580 DGND.n470 DGND.n449 0.0673605
R1581 DGND.n475 DGND.n449 0.0673605
R1582 DGND.n484 DGND.n483 0.0673605
R1583 DGND.n633 DGND.n443 0.0673605
R1584 DGND.n652 DGND.n651 0.0673605
R1585 DGND.n664 DGND.n663 0.0673605
R1586 DGND.n681 DGND.n680 0.0673605
R1587 DGND.n511 DGND.n490 0.0673605
R1588 DGND.n528 DGND.n527 0.0673605
R1589 DGND.n539 DGND.n538 0.0673605
R1590 DGND.n559 DGND.n494 0.0673605
R1591 DGND.n603 DGND.n493 0.0673605
R1592 DGND.n595 DGND.n569 0.0673605
R1593 DGND.n590 DGND.n569 0.0673605
R1594 DGND.n590 DGND.n589 0.0673605
R1595 DGND.n589 DGND.n576 0.0673605
R1596 DGND.n585 DGND.n576 0.0673605
R1597 DGND.n585 DGND.n584 0.0673605
R1598 DGND.n584 DGND.n583 0.0673605
R1599 DGND.n289 DGND.n286 0.0673605
R1600 DGND.n289 DGND.n284 0.0673605
R1601 DGND.n294 DGND.n284 0.0673605
R1602 DGND.n294 DGND.n281 0.0673605
R1603 DGND.n299 DGND.n281 0.0673605
R1604 DGND.n299 DGND.n278 0.0673605
R1605 DGND.n304 DGND.n278 0.0673605
R1606 DGND.n313 DGND.n312 0.0673605
R1607 DGND.n272 DGND.n207 0.0673605
R1608 DGND.n254 DGND.n253 0.0673605
R1609 DGND.n246 DGND.n245 0.0673605
R1610 DGND.n237 DGND.n90 0.0673605
R1611 DGND.n889 DGND.n86 0.0673605
R1612 DGND.n877 DGND.n832 0.0673605
R1613 DGND.n867 DGND.n837 0.0673605
R1614 DGND.n849 DGND.n848 0.0673605
R1615 DGND.n83 DGND.n82 0.0673605
R1616 DGND.n75 DGND.n49 0.0673605
R1617 DGND.n70 DGND.n49 0.0673605
R1618 DGND.n70 DGND.n69 0.0673605
R1619 DGND.n69 DGND.n56 0.0673605
R1620 DGND.n65 DGND.n56 0.0673605
R1621 DGND.n65 DGND.n64 0.0673605
R1622 DGND.n64 DGND.n63 0.0673605
R1623 DGND.n341 DGND.n338 0.0673605
R1624 DGND.n341 DGND.n336 0.0673605
R1625 DGND.n346 DGND.n336 0.0673605
R1626 DGND.n346 DGND.n333 0.0673605
R1627 DGND.n351 DGND.n333 0.0673605
R1628 DGND.n351 DGND.n330 0.0673605
R1629 DGND.n356 DGND.n330 0.0673605
R1630 DGND.n365 DGND.n364 0.0673605
R1631 DGND.n386 DGND.n324 0.0673605
R1632 DGND.n406 DGND.n376 0.0673605
R1633 DGND.n416 DGND.n372 0.0673605
R1634 DGND.n431 DGND.n428 0.0673605
R1635 DGND.n937 DGND.n23 0.0673605
R1636 DGND.n927 DGND.n28 0.0673605
R1637 DGND.n909 DGND.n908 0.0673605
R1638 DGND.n956 DGND.n955 0.0673605
R1639 DGND.n963 DGND.n7 0.0673605
R1640 DGND.n971 DGND.n7 0.0673605
R1641 DGND.n971 DGND.n4 0.0673605
R1642 DGND.n4 DGND.n3 0.0673605
R1643 DGND.n977 DGND.n3 0.0673605
R1644 DGND.n977 DGND.n0 0.0673605
R1645 DGND.n728 DGND.n702 0.0557326
R1646 DGND.n734 DGND.n733 0.0557326
R1647 DGND.n737 DGND.n701 0.0557326
R1648 DGND.n150 DGND.n115 0.0557326
R1649 DGND.n149 DGND.n118 0.0557326
R1650 DGND.n147 DGND.n146 0.0557326
R1651 DGND.n476 DGND.n475 0.0557326
R1652 DGND.n479 DGND.n448 0.0557326
R1653 DGND.n480 DGND.n445 0.0557326
R1654 DGND.n599 DGND.n566 0.0557326
R1655 DGND.n598 DGND.n567 0.0557326
R1656 DGND.n596 DGND.n595 0.0557326
R1657 DGND.n305 DGND.n304 0.0557326
R1658 DGND.n308 DGND.n277 0.0557326
R1659 DGND.n309 DGND.n274 0.0557326
R1660 DGND.n79 DGND.n44 0.0557326
R1661 DGND.n78 DGND.n47 0.0557326
R1662 DGND.n76 DGND.n75 0.0557326
R1663 DGND.n357 DGND.n356 0.0557326
R1664 DGND.n360 DGND.n329 0.0557326
R1665 DGND.n361 DGND.n326 0.0557326
R1666 DGND.n959 DGND.n12 0.0557326
R1667 DGND.n960 DGND.n10 0.0557326
R1668 DGND.n963 DGND.n962 0.0557326
R1669 DGND.n806 DGND.n699 0.0513721
R1670 DGND.n112 DGND.n40 0.0513721
R1671 DGND.n696 DGND.n442 0.0513721
R1672 DGND.n561 DGND.n39 0.0513721
R1673 DGND.n322 DGND.n206 0.0513721
R1674 DGND.n900 DGND.n899 0.0513721
R1675 DGND.n441 DGND.n323 0.0513721
R1676 DGND.n904 DGND.n903 0.0513721
R1677 DGND DGND.n981 0.0499186
R1678 DGND.n686 DGND.n685 0.0484731
R1679 DGND.n614 DGND.n488 0.0484731
R1680 DGND.n818 DGND.n87 0.0484731
R1681 DGND.n819 DGND.n84 0.0484731
R1682 DGND.n775 DGND.n760 0.0470116
R1683 DGND.n773 DGND.n772 0.0470116
R1684 DGND.n764 DGND.n762 0.0470116
R1685 DGND.n769 DGND.n765 0.0470116
R1686 DGND.n199 DGND.n91 0.0470116
R1687 DGND.n198 DGND.n93 0.0470116
R1688 DGND.n195 DGND.n194 0.0470116
R1689 DGND.n192 DGND.n95 0.0470116
R1690 DGND.n667 DGND.n620 0.0470116
R1691 DGND.n668 DGND.n619 0.0470116
R1692 DGND.n677 DGND.n676 0.0470116
R1693 DGND.n679 DGND.n617 0.0470116
R1694 DGND.n518 DGND.n510 0.0470116
R1695 DGND.n519 DGND.n509 0.0470116
R1696 DGND.n524 DGND.n523 0.0470116
R1697 DGND.n526 DGND.n507 0.0470116
R1698 DGND.n244 DGND.n225 0.0470116
R1699 DGND.n242 DGND.n241 0.0470116
R1700 DGND.n229 DGND.n227 0.0470116
R1701 DGND.n238 DGND.n230 0.0470116
R1702 DGND.n885 DGND.n824 0.0470116
R1703 DGND.n884 DGND.n825 0.0470116
R1704 DGND.n881 DGND.n880 0.0470116
R1705 DGND.n878 DGND.n827 0.0470116
R1706 DGND.n417 DGND.n371 0.0470116
R1707 DGND.n420 DGND.n419 0.0470116
R1708 DGND.n423 DGND.n369 0.0470116
R1709 DGND.n424 DGND.n367 0.0470116
R1710 DGND.n17 DGND.n16 0.0470116
R1711 DGND.n945 DGND.n18 0.0470116
R1712 DGND.n944 DGND.n20 0.0470116
R1713 DGND.n941 DGND.n940 0.0470116
R1714 DGND.n938 DGND.n22 0.0470116
R1715 DGND.n739 DGND.n204 0.0441047
R1716 DGND.n807 DGND.n205 0.0441047
R1717 DGND.n799 DGND.n744 0.0441047
R1718 DGND.n798 DGND.n745 0.0441047
R1719 DGND.n795 DGND.n794 0.0441047
R1720 DGND.n790 DGND.n748 0.0441047
R1721 DGND.n789 DGND.n750 0.0441047
R1722 DGND.n176 DGND.n104 0.0441047
R1723 DGND.n175 DGND.n105 0.0441047
R1724 DGND.n171 DGND.n170 0.0441047
R1725 DGND.n167 DGND.n108 0.0441047
R1726 DGND.n166 DGND.n110 0.0441047
R1727 DGND.n158 DGND.n114 0.0441047
R1728 DGND.n157 DGND.n154 0.0441047
R1729 DGND.n485 DGND.n484 0.0441047
R1730 DGND.n692 DGND.n691 0.0441047
R1731 DGND.n636 DGND.n635 0.0441047
R1732 DGND.n639 DGND.n630 0.0441047
R1733 DGND.n640 DGND.n628 0.0441047
R1734 DGND.n647 DGND.n646 0.0441047
R1735 DGND.n650 DGND.n625 0.0441047
R1736 DGND.n544 DGND.n501 0.0441047
R1737 DGND.n545 DGND.n498 0.0441047
R1738 DGND.n550 DGND.n548 0.0441047
R1739 DGND.n549 DGND.n496 0.0441047
R1740 DGND.n555 DGND.n554 0.0441047
R1741 DGND.n492 DGND.n491 0.0441047
R1742 DGND.n604 DGND.n603 0.0441047
R1743 DGND.n314 DGND.n313 0.0441047
R1744 DGND.n318 DGND.n317 0.0441047
R1745 DGND.n268 DGND.n209 0.0441047
R1746 DGND.n267 DGND.n210 0.0441047
R1747 DGND.n264 DGND.n263 0.0441047
R1748 DGND.n259 DGND.n213 0.0441047
R1749 DGND.n258 DGND.n215 0.0441047
R1750 DGND.n862 DGND.n840 0.0441047
R1751 DGND.n861 DGND.n841 0.0441047
R1752 DGND.n857 DGND.n856 0.0441047
R1753 DGND.n853 DGND.n844 0.0441047
R1754 DGND.n852 DGND.n846 0.0441047
R1755 DGND.n896 DGND.n42 0.0441047
R1756 DGND.n895 DGND.n83 0.0441047
R1757 DGND.n366 DGND.n365 0.0441047
R1758 DGND.n437 DGND.n436 0.0441047
R1759 DGND.n388 DGND.n387 0.0441047
R1760 DGND.n393 DGND.n383 0.0441047
R1761 DGND.n392 DGND.n380 0.0441047
R1762 DGND.n379 DGND.n378 0.0441047
R1763 DGND.n399 DGND.n398 0.0441047
R1764 DGND.n922 DGND.n31 0.0441047
R1765 DGND.n921 DGND.n32 0.0441047
R1766 DGND.n917 DGND.n916 0.0441047
R1767 DGND.n913 DGND.n35 0.0441047
R1768 DGND.n912 DGND.n37 0.0441047
R1769 DGND.n15 DGND.n14 0.0441047
R1770 DGND.n955 DGND.n954 0.0441047
R1771 DGND.n783 DGND.n753 0.0353837
R1772 DGND.n781 DGND.n780 0.0353837
R1773 DGND.n777 DGND.n755 0.0353837
R1774 DGND.n182 DGND.n96 0.0353837
R1775 DGND.n100 DGND.n98 0.0353837
R1776 DGND.n186 DGND.n185 0.0353837
R1777 DGND.n658 DGND.n623 0.0353837
R1778 DGND.n659 DGND.n622 0.0353837
R1779 DGND.n663 DGND.n662 0.0353837
R1780 DGND.n681 DGND.n486 0.0353837
R1781 DGND.n686 DGND.n487 0.0353837
R1782 DGND.n610 DGND.n488 0.0353837
R1783 DGND.n609 DGND.n490 0.0353837
R1784 DGND.n528 DGND.n505 0.0353837
R1785 DGND.n535 DGND.n534 0.0353837
R1786 DGND.n537 DGND.n503 0.0353837
R1787 DGND.n252 DGND.n218 0.0353837
R1788 DGND.n250 DGND.n249 0.0353837
R1789 DGND.n246 DGND.n220 0.0353837
R1790 DGND.n814 DGND.n90 0.0353837
R1791 DGND.n815 DGND.n87 0.0353837
R1792 DGND.n85 DGND.n84 0.0353837
R1793 DGND.n890 DGND.n889 0.0353837
R1794 DGND.n868 DGND.n832 0.0353837
R1795 DGND.n836 DGND.n834 0.0353837
R1796 DGND.n872 DGND.n871 0.0353837
R1797 DGND.n408 DGND.n407 0.0353837
R1798 DGND.n412 DGND.n375 0.0353837
R1799 DGND.n411 DGND.n372 0.0353837
R1800 DGND.n928 DGND.n23 0.0353837
R1801 DGND.n27 DGND.n25 0.0353837
R1802 DGND.n932 DGND.n931 0.0353837
R1803 DGND.n804 DGND.n803 0.0324767
R1804 DGND.n784 DGND.n783 0.0324767
R1805 DGND.n781 DGND.n753 0.0324767
R1806 DGND.n780 DGND.n755 0.0324767
R1807 DGND.n182 DGND.n98 0.0324767
R1808 DGND.n186 DGND.n100 0.0324767
R1809 DGND.n185 DGND.n181 0.0324767
R1810 DGND.n162 DGND.n161 0.0324767
R1811 DGND.n695 DGND.n443 0.0324767
R1812 DGND.n652 DGND.n623 0.0324767
R1813 DGND.n659 DGND.n658 0.0324767
R1814 DGND.n662 DGND.n622 0.0324767
R1815 DGND.n487 DGND.n486 0.0324767
R1816 DGND.n610 DGND.n609 0.0324767
R1817 DGND.n534 DGND.n505 0.0324767
R1818 DGND.n535 DGND.n503 0.0324767
R1819 DGND.n538 DGND.n537 0.0324767
R1820 DGND.n560 DGND.n559 0.0324767
R1821 DGND.n321 DGND.n272 0.0324767
R1822 DGND.n253 DGND.n252 0.0324767
R1823 DGND.n250 DGND.n218 0.0324767
R1824 DGND.n249 DGND.n220 0.0324767
R1825 DGND.n815 DGND.n814 0.0324767
R1826 DGND.n890 DGND.n85 0.0324767
R1827 DGND.n868 DGND.n834 0.0324767
R1828 DGND.n872 DGND.n836 0.0324767
R1829 DGND.n871 DGND.n867 0.0324767
R1830 DGND.n848 DGND.n41 0.0324767
R1831 DGND.n440 DGND.n324 0.0324767
R1832 DGND.n408 DGND.n406 0.0324767
R1833 DGND.n407 DGND.n375 0.0324767
R1834 DGND.n412 DGND.n411 0.0324767
R1835 DGND.n928 DGND.n25 0.0324767
R1836 DGND.n932 DGND.n27 0.0324767
R1837 DGND.n931 DGND.n927 0.0324767
R1838 DGND.n908 DGND.n907 0.0324767
R1839 DGND.n205 DGND.n204 0.0237558
R1840 DGND.n807 DGND.n806 0.0237558
R1841 DGND.n744 DGND.n742 0.0237558
R1842 DGND.n799 DGND.n798 0.0237558
R1843 DGND.n795 DGND.n745 0.0237558
R1844 DGND.n794 DGND.n748 0.0237558
R1845 DGND.n790 DGND.n789 0.0237558
R1846 DGND.n785 DGND.n750 0.0237558
R1847 DGND.n104 DGND.n101 0.0237558
R1848 DGND.n176 DGND.n175 0.0237558
R1849 DGND.n171 DGND.n105 0.0237558
R1850 DGND.n170 DGND.n108 0.0237558
R1851 DGND.n167 DGND.n166 0.0237558
R1852 DGND.n163 DGND.n110 0.0237558
R1853 DGND.n114 DGND.n112 0.0237558
R1854 DGND.n158 DGND.n157 0.0237558
R1855 DGND.n692 DGND.n485 0.0237558
R1856 DGND.n691 DGND.n442 0.0237558
R1857 DGND.n635 DGND.n633 0.0237558
R1858 DGND.n636 DGND.n630 0.0237558
R1859 DGND.n640 DGND.n639 0.0237558
R1860 DGND.n646 DGND.n628 0.0237558
R1861 DGND.n647 DGND.n625 0.0237558
R1862 DGND.n651 DGND.n650 0.0237558
R1863 DGND.n539 DGND.n501 0.0237558
R1864 DGND.n545 DGND.n544 0.0237558
R1865 DGND.n548 DGND.n498 0.0237558
R1866 DGND.n550 DGND.n549 0.0237558
R1867 DGND.n555 DGND.n496 0.0237558
R1868 DGND.n554 DGND.n494 0.0237558
R1869 DGND.n561 DGND.n491 0.0237558
R1870 DGND.n604 DGND.n492 0.0237558
R1871 DGND.n318 DGND.n314 0.0237558
R1872 DGND.n317 DGND.n206 0.0237558
R1873 DGND.n209 DGND.n207 0.0237558
R1874 DGND.n268 DGND.n267 0.0237558
R1875 DGND.n264 DGND.n210 0.0237558
R1876 DGND.n263 DGND.n213 0.0237558
R1877 DGND.n259 DGND.n258 0.0237558
R1878 DGND.n254 DGND.n215 0.0237558
R1879 DGND.n840 DGND.n837 0.0237558
R1880 DGND.n862 DGND.n861 0.0237558
R1881 DGND.n857 DGND.n841 0.0237558
R1882 DGND.n856 DGND.n844 0.0237558
R1883 DGND.n853 DGND.n852 0.0237558
R1884 DGND.n849 DGND.n846 0.0237558
R1885 DGND.n899 DGND.n42 0.0237558
R1886 DGND.n896 DGND.n895 0.0237558
R1887 DGND.n437 DGND.n366 0.0237558
R1888 DGND.n436 DGND.n323 0.0237558
R1889 DGND.n388 DGND.n386 0.0237558
R1890 DGND.n387 DGND.n383 0.0237558
R1891 DGND.n393 DGND.n392 0.0237558
R1892 DGND.n380 DGND.n379 0.0237558
R1893 DGND.n399 DGND.n378 0.0237558
R1894 DGND.n398 DGND.n376 0.0237558
R1895 DGND.n31 DGND.n28 0.0237558
R1896 DGND.n922 DGND.n921 0.0237558
R1897 DGND.n917 DGND.n32 0.0237558
R1898 DGND.n916 DGND.n35 0.0237558
R1899 DGND.n913 DGND.n912 0.0237558
R1900 DGND.n909 DGND.n37 0.0237558
R1901 DGND.n904 DGND.n15 0.0237558
R1902 DGND.n954 DGND.n14 0.0237558
R1903 DGND.n776 DGND.n775 0.0208488
R1904 DGND.n773 DGND.n760 0.0208488
R1905 DGND.n772 DGND.n762 0.0208488
R1906 DGND.n765 DGND.n764 0.0208488
R1907 DGND.n769 DGND.n768 0.0208488
R1908 DGND.n202 DGND.n91 0.0208488
R1909 DGND.n199 DGND.n198 0.0208488
R1910 DGND.n195 DGND.n93 0.0208488
R1911 DGND.n194 DGND.n95 0.0208488
R1912 DGND.n192 DGND.n191 0.0208488
R1913 DGND.n664 DGND.n620 0.0208488
R1914 DGND.n668 DGND.n667 0.0208488
R1915 DGND.n676 DGND.n619 0.0208488
R1916 DGND.n677 DGND.n617 0.0208488
R1917 DGND.n680 DGND.n679 0.0208488
R1918 DGND.n511 DGND.n510 0.0208488
R1919 DGND.n519 DGND.n518 0.0208488
R1920 DGND.n523 DGND.n509 0.0208488
R1921 DGND.n524 DGND.n507 0.0208488
R1922 DGND.n527 DGND.n526 0.0208488
R1923 DGND.n245 DGND.n244 0.0208488
R1924 DGND.n242 DGND.n225 0.0208488
R1925 DGND.n241 DGND.n227 0.0208488
R1926 DGND.n230 DGND.n229 0.0208488
R1927 DGND.n238 DGND.n237 0.0208488
R1928 DGND.n824 DGND.n86 0.0208488
R1929 DGND.n885 DGND.n884 0.0208488
R1930 DGND.n881 DGND.n825 0.0208488
R1931 DGND.n880 DGND.n827 0.0208488
R1932 DGND.n878 DGND.n877 0.0208488
R1933 DGND.n417 DGND.n416 0.0208488
R1934 DGND.n419 DGND.n371 0.0208488
R1935 DGND.n420 DGND.n369 0.0208488
R1936 DGND.n424 DGND.n423 0.0208488
R1937 DGND.n427 DGND.n367 0.0208488
R1938 DGND.n428 DGND.n16 0.0208488
R1939 DGND.n949 DGND.n17 0.0208488
R1940 DGND.n948 DGND.n18 0.0208488
R1941 DGND.n945 DGND.n944 0.0208488
R1942 DGND.n941 DGND.n20 0.0208488
R1943 DGND.n940 DGND.n22 0.0208488
R1944 DGND.n938 DGND.n937 0.0208488
R1945 DGND DGND.n0 0.0179419
R1946 DGND.n804 DGND.n699 0.0164884
R1947 DGND.n161 DGND.n40 0.0164884
R1948 DGND.n696 DGND.n695 0.0164884
R1949 DGND.n560 DGND.n39 0.0164884
R1950 DGND.n322 DGND.n321 0.0164884
R1951 DGND.n900 DGND.n41 0.0164884
R1952 DGND.n441 DGND.n440 0.0164884
R1953 DGND.n907 DGND.n903 0.0164884
R1954 DGND.n733 DGND.n702 0.0121279
R1955 DGND.n734 DGND.n701 0.0121279
R1956 DGND.n738 DGND.n737 0.0121279
R1957 DGND.n153 DGND.n115 0.0121279
R1958 DGND.n150 DGND.n149 0.0121279
R1959 DGND.n147 DGND.n118 0.0121279
R1960 DGND.n476 DGND.n448 0.0121279
R1961 DGND.n480 DGND.n479 0.0121279
R1962 DGND.n483 DGND.n445 0.0121279
R1963 DGND.n566 DGND.n493 0.0121279
R1964 DGND.n599 DGND.n598 0.0121279
R1965 DGND.n596 DGND.n567 0.0121279
R1966 DGND.n305 DGND.n277 0.0121279
R1967 DGND.n309 DGND.n308 0.0121279
R1968 DGND.n312 DGND.n274 0.0121279
R1969 DGND.n82 DGND.n44 0.0121279
R1970 DGND.n79 DGND.n78 0.0121279
R1971 DGND.n76 DGND.n47 0.0121279
R1972 DGND.n357 DGND.n329 0.0121279
R1973 DGND.n361 DGND.n360 0.0121279
R1974 DGND.n364 DGND.n326 0.0121279
R1975 DGND.n956 DGND.n12 0.0121279
R1976 DGND.n960 DGND.n959 0.0121279
R1977 DGND.n962 DGND.n10 0.0121279
R1978 DVDD.n877 DVDD.t419 1255.17
R1979 DVDD.n876 DVDD.t33 1255.17
R1980 DVDD.t428 DVDD.t432 1198.6
R1981 DVDD.t174 DVDD.t8 1198.6
R1982 DVDD.n802 DVDD.t302 1090.58
R1983 DVDD.t263 DVDD.t192 1038.79
R1984 DVDD.t146 DVDD.t461 1038.79
R1985 DVDD.t242 DVDD.t67 944.082
R1986 DVDD.t7 DVDD.t263 944.082
R1987 DVDD.t461 DVDD.t60 944.082
R1988 DVDD.t24 DVDD.t519 944.082
R1989 DVDD.n334 DVDD.t242 896.73
R1990 DVDD.n333 DVDD.t24 896.73
R1991 DVDD.n326 DVDD.t482 842.073
R1992 DVDD.n734 DVDD.t368 842.073
R1993 DVDD.n151 DVDD.t362 842.073
R1994 DVDD.n79 DVDD.t518 842.073
R1995 DVDD.n42 DVDD.t293 842.073
R1996 DVDD.n719 DVDD.t409 842.073
R1997 DVDD.n648 DVDD.t205 842.073
R1998 DVDD.n508 DVDD.t77 842.073
R1999 DVDD.n586 DVDD.t489 842.073
R2000 DVDD.n470 DVDD.t387 842.073
R2001 DVDD.n401 DVDD.t385 842.073
R2002 DVDD.n193 DVDD.t523 842.073
R2003 DVDD.n350 DVDD.t307 842.073
R2004 DVDD.n268 DVDD.t59 842.073
R2005 DVDD.n286 DVDD.t299 842.073
R2006 DVDD.n264 DVDD.t82 842.073
R2007 DVDD.n334 DVDD.t358 799.066
R2008 DVDD.t376 DVDD.n333 799.066
R2009 DVDD.t377 DVDD.t119 781.308
R2010 DVDD.t326 DVDD.t51 781.308
R2011 DVDD.t300 DVDD.n442 737.275
R2012 DVDD.n378 DVDD.t508 737.275
R2013 DVDD.n729 DVDD.t318 703.981
R2014 DVDD.n149 DVDD.t74 703.981
R2015 DVDD.n73 DVDD.t229 703.981
R2016 DVDD.n36 DVDD.t471 703.981
R2017 DVDD.n724 DVDD.t521 703.981
R2018 DVDD.n646 DVDD.t207 703.981
R2019 DVDD.n564 DVDD.t403 703.981
R2020 DVDD.n581 DVDD.t30 703.981
R2021 DVDD.n475 DVDD.t64 703.981
R2022 DVDD.n399 DVDD.t389 703.981
R2023 DVDD.n248 DVDD.t278 703.981
R2024 DVDD.n345 DVDD.t139 703.981
R2025 DVDD.n922 DVDD.t95 703.981
R2026 DVDD.n899 DVDD.t429 703.981
R2027 DVDD.n854 DVDD.t175 703.981
R2028 DVDD.n831 DVDD.t309 703.981
R2029 DVDD.n757 DVDD.t39 697.465
R2030 DVDD.n793 DVDD.t337 697.465
R2031 DVDD.n116 DVDD.t41 697.465
R2032 DVDD.n76 DVDD.t345 697.465
R2033 DVDD.n491 DVDD.t437 697.465
R2034 DVDD.n682 DVDD.t55 697.465
R2035 DVDD.n530 DVDD.t360 697.465
R2036 DVDD.n609 DVDD.t66 697.465
R2037 DVDD.n184 DVDD.t464 697.465
R2038 DVDD.n436 DVDD.t90 697.465
R2039 DVDD.n215 DVDD.t286 697.465
R2040 DVDD.n373 DVDD.t99 697.465
R2041 DVDD.n901 DVDD.t433 697.465
R2042 DVDD.n879 DVDD.t420 697.465
R2043 DVDD.n874 DVDD.t34 697.465
R2044 DVDD.n851 DVDD.t9 697.465
R2045 DVDD.n741 DVDD.t364 663.062
R2046 DVDD.n142 DVDD.t383 663.062
R2047 DVDD.n65 DVDD.t164 663.062
R2048 DVDD.n816 DVDD.t534 663.062
R2049 DVDD.n485 DVDD.t158 663.062
R2050 DVDD.n639 DVDD.t181 663.062
R2051 DVDD.n548 DVDD.t513 663.062
R2052 DVDD.n572 DVDD.t236 663.062
R2053 DVDD.n178 DVDD.t416 663.062
R2054 DVDD.n392 DVDD.t414 663.062
R2055 DVDD.n232 DVDD.t439 663.062
R2056 DVDD.n256 DVDD.t15 663.062
R2057 DVDD.n912 DVDD.t71 663.062
R2058 DVDD.n12 DVDD.t478 663.062
R2059 DVDD.n21 DVDD.t209 663.062
R2060 DVDD.n30 DVDD.t156 663.062
R2061 DVDD.t162 DVDD.t46 633.333
R2062 DVDD.t220 DVDD.t457 633.333
R2063 DVDD.n632 DVDD.n631 629.801
R2064 DVDD.n534 DVDD.n523 629.801
R2065 DVDD.n272 DVDD.n271 629.801
R2066 DVDD.n282 DVDD.n281 629.801
R2067 DVDD.n161 DVDD.n160 598.965
R2068 DVDD.n156 DVDD.n155 598.965
R2069 DVDD.n774 DVDD.n773 598.965
R2070 DVDD.n783 DVDD.n782 598.965
R2071 DVDD.n105 DVDD.n64 598.965
R2072 DVDD.n94 DVDD.n67 598.965
R2073 DVDD.n49 DVDD.n48 598.965
R2074 DVDD.n47 DVDD.n45 598.965
R2075 DVDD.n713 DVDD.n484 598.965
R2076 DVDD.n706 DVDD.n488 598.965
R2077 DVDD.n664 DVDD.n663 598.965
R2078 DVDD.n673 DVDD.n672 598.965
R2079 DVDD.n516 DVDD.n515 598.965
R2080 DVDD.n513 DVDD.n512 598.965
R2081 DVDD.n599 DVDD.n571 598.965
R2082 DVDD.n592 DVDD.n577 598.965
R2083 DVDD.n464 DVDD.n177 598.965
R2084 DVDD.n457 DVDD.n181 598.965
R2085 DVDD.n417 DVDD.n416 598.965
R2086 DVDD.n426 DVDD.n425 598.965
R2087 DVDD.n201 DVDD.n200 598.965
R2088 DVDD.n198 DVDD.n197 598.965
R2089 DVDD.n363 DVDD.n255 598.965
R2090 DVDD.n356 DVDD.n261 598.965
R2091 DVDD.n915 DVDD.n914 598.965
R2092 DVDD.n5 DVDD.n4 598.965
R2093 DVDD.n892 DVDD.n11 598.965
R2094 DVDD.n886 DVDD.n14 598.965
R2095 DVDD.n867 DVDD.n20 598.965
R2096 DVDD.n861 DVDD.n23 598.965
R2097 DVDD.n844 DVDD.n29 598.965
R2098 DVDD.n838 DVDD.n32 598.965
R2099 DVDD.t81 DVDD.t257 556.386
R2100 DVDD.t358 DVDD.t298 556.386
R2101 DVDD.t58 DVDD.t376 556.386
R2102 DVDD.t481 DVDD.t491 556.386
R2103 DVDD.t477 DVDD.t369 556.386
R2104 DVDD.t70 DVDD.t68 556.386
R2105 DVDD.t155 DVDD.t16 556.386
R2106 DVDD.t208 DVDD.t244 556.386
R2107 DVDD.t128 DVDD.n802 497.197
R2108 DVDD.n801 DVDD.t444 346.262
R2109 DVDD.n788 DVDD.t320 340.301
R2110 DVDD.n110 DVDD.t451 340.301
R2111 DVDD.n431 DVDD.t469 340.301
R2112 DVDD.n208 DVDD.t199 340.301
R2113 DVDD.t38 DVDD.t186 338.863
R2114 DVDD.t344 DVDD.t137 338.863
R2115 DVDD.t436 DVDD.t434 338.863
R2116 DVDD.t136 DVDD.t65 338.863
R2117 DVDD.t463 DVDD.t222 338.863
R2118 DVDD.t490 DVDD.t98 338.863
R2119 DVDD.n324 DVDD.n323 324.74
R2120 DVDD.n166 DVDD.n165 324.74
R2121 DVDD.n768 DVDD.n146 324.74
R2122 DVDD.n89 DVDD.n70 324.74
R2123 DVDD.n821 DVDD.n43 324.74
R2124 DVDD.n482 DVDD.n481 324.74
R2125 DVDD.n658 DVDD.n643 324.74
R2126 DVDD.n510 DVDD.n509 324.74
R2127 DVDD.n575 DVDD.n574 324.74
R2128 DVDD.n175 DVDD.n174 324.74
R2129 DVDD.n411 DVDD.n396 324.74
R2130 DVDD.n195 DVDD.n194 324.74
R2131 DVDD.n259 DVDD.n258 324.74
R2132 DVDD.n318 DVDD.n270 324.74
R2133 DVDD.n284 DVDD.n283 324.74
R2134 DVDD.n338 DVDD.n266 324.74
R2135 DVDD.t190 DVDD.t326 322.587
R2136 DVDD.t51 DVDD.t148 322.587
R2137 DVDD.n131 DVDD.n130 320.976
R2138 DVDD.n58 DVDD.n57 320.976
R2139 DVDD.n381 DVDD.n380 320.976
R2140 DVDD.n210 DVDD.n209 320.976
R2141 DVDD.t43 DVDD.t390 316.668
R2142 DVDD.t479 DVDD.t297 316.668
R2143 DVDD.t46 DVDD.t190 304.829
R2144 DVDD.t148 DVDD.t220 304.829
R2145 DVDD.t192 DVDD.t230 284.113
R2146 DVDD.t4 DVDD.t146 284.113
R2147 DVDD.t419 DVDD.t291 284.113
R2148 DVDD.t144 DVDD.t240 284.113
R2149 DVDD.t432 DVDD.t405 284.113
R2150 DVDD.t480 DVDD.t80 284.113
R2151 DVDD.t150 DVDD.t346 284.113
R2152 DVDD.t8 DVDD.t123 284.113
R2153 DVDD.t265 DVDD.t349 284.113
R2154 DVDD.t33 DVDD.t467 284.113
R2155 DVDD.t324 DVDD.t382 278.193
R2156 DVDD.t178 DVDD.t163 278.193
R2157 DVDD.t294 DVDD.t180 278.193
R2158 DVDD.t512 DVDD.t524 278.193
R2159 DVDD.t338 DVDD.t413 278.193
R2160 DVDD.t438 DVDD.t453 278.193
R2161 DVDD.t535 DVDD.t428 266.356
R2162 DVDD.t404 DVDD.t94 266.356
R2163 DVDD.t248 DVDD.t308 266.356
R2164 DVDD.t75 DVDD.t174 266.356
R2165 DVDD.n331 DVDD.t25 264.812
R2166 DVDD.n316 DVDD.t462 264.812
R2167 DVDD.n291 DVDD.t264 264.812
R2168 DVDD.n336 DVDD.t243 264.812
R2169 DVDD.t240 DVDD.t426 263.397
R2170 DVDD.t80 DVDD.t430 263.397
R2171 DVDD.t346 DVDD.t310 263.397
R2172 DVDD.t349 DVDD.t504 263.397
R2173 DVDD.t186 DVDD.t73 260.437
R2174 DVDD.t137 DVDD.t228 260.437
R2175 DVDD.t434 DVDD.t206 260.437
R2176 DVDD.t402 DVDD.t136 260.437
R2177 DVDD.t222 DVDD.t388 260.437
R2178 DVDD.t277 DVDD.t490 260.437
R2179 DVDD.n158 DVDD.t79 255.904
R2180 DVDD.n140 DVDD.t239 255.904
R2181 DVDD.n124 DVDD.t303 255.904
R2182 DVDD.n100 DVDD.t351 255.904
R2183 DVDD.n51 DVDD.t348 255.904
R2184 DVDD.n701 DVDD.t374 255.904
R2185 DVDD.n637 DVDD.t397 255.904
R2186 DVDD.n543 DVDD.t112 255.904
R2187 DVDD.n603 DVDD.t530 255.904
R2188 DVDD.n452 DVDD.t315 255.904
R2189 DVDD.n390 DVDD.t216 255.904
R2190 DVDD.n227 DVDD.t322 255.904
R2191 DVDD.n367 DVDD.t196 255.904
R2192 DVDD.n797 DVDD.t445 249.362
R2193 DVDD.n120 DVDD.t129 249.362
R2194 DVDD.n440 DVDD.t301 249.362
R2195 DVDD.n211 DVDD.t509 249.362
R2196 DVDD.t44 DVDD.t81 248.599
R2197 DVDD.t273 DVDD.t44 248.599
R2198 DVDD.t67 DVDD.t273 248.599
R2199 DVDD.t298 DVDD.t281 248.599
R2200 DVDD.t281 DVDD.t279 248.599
R2201 DVDD.t279 DVDD.t7 248.599
R2202 DVDD.t60 DVDD.t87 248.599
R2203 DVDD.t87 DVDD.t91 248.599
R2204 DVDD.t91 DVDD.t58 248.599
R2205 DVDD.t519 DVDD.t121 248.599
R2206 DVDD.t121 DVDD.t100 248.599
R2207 DVDD.t100 DVDD.t481 248.599
R2208 DVDD.t426 DVDD.t142 248.599
R2209 DVDD.t142 DVDD.t477 248.599
R2210 DVDD.t369 DVDD.t421 248.599
R2211 DVDD.t421 DVDD.t145 248.599
R2212 DVDD.t145 DVDD.t535 248.599
R2213 DVDD.t430 DVDD.t497 248.599
R2214 DVDD.t497 DVDD.t70 248.599
R2215 DVDD.t68 DVDD.t536 248.599
R2216 DVDD.t536 DVDD.t496 248.599
R2217 DVDD.t496 DVDD.t404 248.599
R2218 DVDD.t410 DVDD.t248 248.599
R2219 DVDD.t160 DVDD.t410 248.599
R2220 DVDD.t16 DVDD.t160 248.599
R2221 DVDD.t379 DVDD.t155 248.599
R2222 DVDD.t310 DVDD.t379 248.599
R2223 DVDD.t268 DVDD.t75 248.599
R2224 DVDD.t35 DVDD.t268 248.599
R2225 DVDD.t244 DVDD.t35 248.599
R2226 DVDD.t266 DVDD.t208 248.599
R2227 DVDD.t504 DVDD.t266 248.599
R2228 DVDD.n802 DVDD.n122 240.078
R2229 DVDD.n333 DVDD.n332 240.065
R2230 DVDD.n335 DVDD.n334 240.065
R2231 DVDD.n497 DVDD.n496 235.248
R2232 DVDD.n620 DVDD.n499 235.248
R2233 DVDD.n305 DVDD.n276 235.248
R2234 DVDD.n302 DVDD.n278 235.248
R2235 DVDD.n753 DVDD.n752 226.786
R2236 DVDD.n801 DVDD.n800 226.786
R2237 DVDD.n804 DVDD.n803 226.786
R2238 DVDD.n613 DVDD.n612 226.786
R2239 DVDD.n693 DVDD.n692 226.786
R2240 DVDD.n691 DVDD.n690 226.786
R2241 DVDD.n615 DVDD.n614 226.786
R2242 DVDD.n444 DVDD.n443 226.786
R2243 DVDD.n377 DVDD.n376 226.786
R2244 DVDD.t230 DVDD.t162 213.084
R2245 DVDD.t457 DVDD.t4 213.084
R2246 DVDD.t291 DVDD.t144 213.084
R2247 DVDD.t405 DVDD.t480 213.084
R2248 DVDD.t123 DVDD.t150 213.084
R2249 DVDD.t467 DVDD.t265 213.084
R2250 DVDD.t363 DVDD.t6 210.125
R2251 DVDD.t533 DVDD.t18 210.125
R2252 DVDD.t157 DVDD.t381 210.125
R2253 DVDD.t235 DVDD.t53 210.125
R2254 DVDD.t415 DVDD.t159 210.125
R2255 DVDD.t14 DVDD.t93 210.125
R2256 DVDD.t119 DVDD.t356 159.321
R2257 DVDD.t446 DVDD.t377 159.321
R2258 DVDD.t398 DVDD.t251 142.056
R2259 DVDD.t3 DVDD.t375 142.056
R2260 DVDD.t203 DVDD.t528 142.056
R2261 DVDD.t110 DVDD.t127 142.056
R2262 DVDD.t214 DVDD.t130 142.056
R2263 DVDD.t221 DVDD.t316 142.056
R2264 DVDD.t47 DVDD.t194 142.056
R2265 DVDD.t258 DVDD.t323 142.056
R2266 DVDD.t460 DVDD.t22 142.056
R2267 DVDD.t213 DVDD.t26 142.056
R2268 DVDD.t269 DVDD.t241 142.056
R2269 DVDD.t484 DVDD.t262 142.056
R2270 DVDD.t435 DVDD.t317 133.179
R2271 DVDD.t532 DVDD.t470 133.179
R2272 DVDD.t423 DVDD.t520 133.179
R2273 DVDD.t312 DVDD.t29 133.179
R2274 DVDD.t13 DVDD.t63 133.179
R2275 DVDD.t335 DVDD.t138 133.179
R2276 DVDD.t151 DVDD.t398 131.698
R2277 DVDD.t255 DVDD.t110 131.698
R2278 DVDD.t333 DVDD.t214 131.698
R2279 DVDD.t323 DVDD.t331 131.698
R2280 DVDD.t442 DVDD.t460 131.698
R2281 DVDD.t262 DVDD.t275 131.698
R2282 DVDD.t304 DVDD.t444 124.299
R2283 DVDD.t252 DVDD.t151 124.299
R2284 DVDD.t106 DVDD.t1 124.299
R2285 DVDD.t1 DVDD.t363 124.299
R2286 DVDD.t200 DVDD.t533 124.299
R2287 DVDD.t492 DVDD.t200 124.299
R2288 DVDD.t124 DVDD.t255 124.299
R2289 DVDD.t249 DVDD.t128 124.299
R2290 DVDD.t132 DVDD.t333 124.299
R2291 DVDD.t499 DVDD.t218 124.299
R2292 DVDD.t218 DVDD.t157 124.299
R2293 DVDD.t48 DVDD.t235 124.299
R2294 DVDD.t10 DVDD.t48 124.299
R2295 DVDD.t331 DVDD.t259 124.299
R2296 DVDD.t455 DVDD.t300 124.299
R2297 DVDD.t20 DVDD.t442 124.299
R2298 DVDD.t61 DVDD.t211 124.299
R2299 DVDD.t211 DVDD.t415 124.299
R2300 DVDD.t270 DVDD.t14 124.299
R2301 DVDD.t140 DVDD.t270 124.299
R2302 DVDD.t275 DVDD.t485 124.299
R2303 DVDD.t508 DVDD.t223 124.299
R2304 DVDD.n496 DVDD.t357 123.507
R2305 DVDD.n499 DVDD.t447 123.507
R2306 DVDD.n276 DVDD.t149 123.507
R2307 DVDD.n278 DVDD.t191 123.507
R2308 DVDD.t375 DVDD.t78 118.38
R2309 DVDD.t528 DVDD.t347 118.38
R2310 DVDD.t316 DVDD.t373 118.38
R2311 DVDD.t194 DVDD.t529 118.38
R2312 DVDD.t26 DVDD.t314 118.38
R2313 DVDD.t241 DVDD.t195 118.38
R2314 DVDD.t225 DVDD.t324 115.421
R2315 DVDD.t417 DVDD.t176 115.421
R2316 DVDD.t424 DVDD.t254 115.421
R2317 DVDD.t361 DVDD.t165 115.421
R2318 DVDD.t517 DVDD.t247 115.421
R2319 DVDD.t83 DVDD.t126 115.421
R2320 DVDD.t153 DVDD.t474 115.421
R2321 DVDD.t501 DVDD.t178 115.421
R2322 DVDD.t390 DVDD.n691 115.421
R2323 DVDD.t476 DVDD.t294 115.421
R2324 DVDD.t85 DVDD.t113 115.421
R2325 DVDD.t104 DVDD.t131 115.421
R2326 DVDD.t204 DVDD.t19 115.421
R2327 DVDD.t290 DVDD.t76 115.421
R2328 DVDD.t261 DVDD.t340 115.421
R2329 DVDD.t56 DVDD.t226 115.421
R2330 DVDD.t524 DVDD.t237 115.421
R2331 DVDD.n614 DVDD.t479 115.421
R2332 DVDD.t289 DVDD.t338 115.421
R2333 DVDD.t371 DVDD.t440 115.421
R2334 DVDD.t31 DVDD.t23 115.421
R2335 DVDD.t384 DVDD.t401 115.421
R2336 DVDD.t452 DVDD.t522 115.421
R2337 DVDD.t487 DVDD.t172 115.421
R2338 DVDD.t283 DVDD.t342 115.421
R2339 DVDD.t453 DVDD.t514 115.421
R2340 DVDD.t302 DVDD.n801 113.942
R2341 DVDD.t296 DVDD.t352 110.981
R2342 DVDD.t510 DVDD.t328 110.981
R2343 DVDD.t12 DVDD.t3 106.543
R2344 DVDD.t232 DVDD.t203 106.543
R2345 DVDD.t406 DVDD.t221 106.543
R2346 DVDD.t72 DVDD.t47 106.543
R2347 DVDD.t483 DVDD.t213 106.543
R2348 DVDD.t246 DVDD.t269 106.543
R2349 DVDD.t134 DVDD.t336 87.3058
R2350 DVDD.t319 DVDD.t187 87.3058
R2351 DVDD.t450 DVDD.t393 87.3058
R2352 DVDD.t399 DVDD.t40 87.3058
R2353 DVDD.t506 DVDD.t89 87.3058
R2354 DVDD.t468 DVDD.t197 87.3058
R2355 DVDD.t37 DVDD.t198 87.3058
R2356 DVDD.t285 DVDD.t526 87.3058
R2357 DVDD.n631 DVDD.t353 86.7743
R2358 DVDD.n523 DVDD.t511 86.7743
R2359 DVDD.n271 DVDD.t5 86.7743
R2360 DVDD.n281 DVDD.t231 86.7743
R2361 DVDD.n752 DVDD.t12 81.3868
R2362 DVDD.n803 DVDD.t232 81.3868
R2363 DVDD.n692 DVDD.t406 81.3868
R2364 DVDD.n613 DVDD.t72 81.3868
R2365 DVDD.n443 DVDD.t483 81.3868
R2366 DVDD.n377 DVDD.t246 81.3868
R2367 DVDD.t382 DVDD.t238 78.4273
R2368 DVDD.t163 DVDD.t350 78.4273
R2369 DVDD.t180 DVDD.t396 78.4273
R2370 DVDD.t111 DVDD.t512 78.4273
R2371 DVDD.t413 DVDD.t215 78.4273
R2372 DVDD.t321 DVDD.t438 78.4273
R2373 DVDD.t317 DVDD.t531 76.9475
R2374 DVDD.t470 DVDD.t171 76.9475
R2375 DVDD.t520 DVDD.t42 76.9475
R2376 DVDD.t29 DVDD.t170 76.9475
R2377 DVDD.t63 DVDD.t313 76.9475
R2378 DVDD.t138 DVDD.t407 76.9475
R2379 DVDD.t54 DVDD.t43 75.4678
R2380 DVDD.t130 DVDD.t354 75.4678
R2381 DVDD.t448 DVDD.t258 75.4678
R2382 DVDD.t297 DVDD.t359 75.4678
R2383 DVDD.t6 DVDD.t117 68.069
R2384 DVDD.t96 DVDD.t458 68.069
R2385 DVDD.t287 DVDD.t0 68.069
R2386 DVDD.t367 DVDD.t435 68.069
R2387 DVDD.t292 DVDD.t532 68.069
R2388 DVDD.t394 DVDD.t202 68.069
R2389 DVDD.t411 DVDD.t494 68.069
R2390 DVDD.t18 DVDD.t329 68.069
R2391 DVDD.t381 DVDD.t182 68.069
R2392 DVDD.t184 DVDD.t465 68.069
R2393 DVDD.t108 DVDD.t217 68.069
R2394 DVDD.t408 DVDD.t423 68.069
R2395 DVDD.t488 DVDD.t312 68.069
R2396 DVDD.t472 DVDD.t50 68.069
R2397 DVDD.t391 DVDD.t168 68.069
R2398 DVDD.t53 DVDD.t233 68.069
R2399 DVDD.t159 DVDD.t365 68.069
R2400 DVDD.t115 DVDD.t102 68.069
R2401 DVDD.t188 DVDD.t210 68.069
R2402 DVDD.t386 DVDD.t13 68.069
R2403 DVDD.t306 DVDD.t335 68.069
R2404 DVDD.t27 DVDD.t272 68.069
R2405 DVDD.t166 DVDD.t515 68.069
R2406 DVDD.t93 DVDD.t502 68.069
R2407 DVDD.n631 DVDD.t355 68.0124
R2408 DVDD.n523 DVDD.t449 68.0124
R2409 DVDD.n271 DVDD.t147 68.0124
R2410 DVDD.n281 DVDD.t193 68.0124
R2411 DVDD.n160 DVDD.t118 63.3219
R2412 DVDD.n160 DVDD.t459 63.3219
R2413 DVDD.n155 DVDD.t107 63.3219
R2414 DVDD.n155 DVDD.t2 63.3219
R2415 DVDD.n773 DVDD.t325 63.3219
R2416 DVDD.n773 DVDD.t177 63.3219
R2417 DVDD.n782 DVDD.t152 63.3219
R2418 DVDD.n782 DVDD.t253 63.3219
R2419 DVDD.n64 DVDD.t125 63.3219
R2420 DVDD.n64 DVDD.t256 63.3219
R2421 DVDD.n67 DVDD.t475 63.3219
R2422 DVDD.n67 DVDD.t179 63.3219
R2423 DVDD.n48 DVDD.t201 63.3219
R2424 DVDD.n48 DVDD.t493 63.3219
R2425 DVDD.n45 DVDD.t495 63.3219
R2426 DVDD.n45 DVDD.t330 63.3219
R2427 DVDD.n484 DVDD.t183 63.3219
R2428 DVDD.n484 DVDD.t466 63.3219
R2429 DVDD.n488 DVDD.t500 63.3219
R2430 DVDD.n488 DVDD.t219 63.3219
R2431 DVDD.n663 DVDD.t295 63.3219
R2432 DVDD.n663 DVDD.t114 63.3219
R2433 DVDD.n672 DVDD.t334 63.3219
R2434 DVDD.n672 DVDD.t133 63.3219
R2435 DVDD.n515 DVDD.t260 63.3219
R2436 DVDD.n515 DVDD.t332 63.3219
R2437 DVDD.n512 DVDD.t57 63.3219
R2438 DVDD.n512 DVDD.t525 63.3219
R2439 DVDD.n571 DVDD.t49 63.3219
R2440 DVDD.n571 DVDD.t11 63.3219
R2441 DVDD.n577 DVDD.t169 63.3219
R2442 DVDD.n577 DVDD.t234 63.3219
R2443 DVDD.n177 DVDD.t366 63.3219
R2444 DVDD.n177 DVDD.t103 63.3219
R2445 DVDD.n181 DVDD.t62 63.3219
R2446 DVDD.n181 DVDD.t212 63.3219
R2447 DVDD.n416 DVDD.t339 63.3219
R2448 DVDD.n416 DVDD.t441 63.3219
R2449 DVDD.n425 DVDD.t443 63.3219
R2450 DVDD.n425 DVDD.t21 63.3219
R2451 DVDD.n200 DVDD.t486 63.3219
R2452 DVDD.n200 DVDD.t276 63.3219
R2453 DVDD.n197 DVDD.t284 63.3219
R2454 DVDD.n197 DVDD.t454 63.3219
R2455 DVDD.n255 DVDD.t271 63.3219
R2456 DVDD.n255 DVDD.t141 63.3219
R2457 DVDD.n261 DVDD.t516 63.3219
R2458 DVDD.n261 DVDD.t503 63.3219
R2459 DVDD.n914 DVDD.t69 63.3219
R2460 DVDD.n914 DVDD.t537 63.3219
R2461 DVDD.n4 DVDD.t431 63.3219
R2462 DVDD.n4 DVDD.t498 63.3219
R2463 DVDD.n11 DVDD.t370 63.3219
R2464 DVDD.n11 DVDD.t422 63.3219
R2465 DVDD.n14 DVDD.t427 63.3219
R2466 DVDD.n14 DVDD.t143 63.3219
R2467 DVDD.n20 DVDD.t267 63.3219
R2468 DVDD.n20 DVDD.t505 63.3219
R2469 DVDD.n23 DVDD.t36 63.3219
R2470 DVDD.n23 DVDD.t245 63.3219
R2471 DVDD.n29 DVDD.t380 63.3219
R2472 DVDD.n29 DVDD.t311 63.3219
R2473 DVDD.n32 DVDD.t161 63.3219
R2474 DVDD.n32 DVDD.t17 63.3219
R2475 DVDD.n752 DVDD.t38 60.6703
R2476 DVDD.n803 DVDD.t344 60.6703
R2477 DVDD.n692 DVDD.t436 60.6703
R2478 DVDD.t65 DVDD.n613 60.6703
R2479 DVDD.n443 DVDD.t463 60.6703
R2480 DVDD.t98 DVDD.n377 60.6703
R2481 DVDD.t117 DVDD.t96 56.231
R2482 DVDD.t458 DVDD.t287 56.231
R2483 DVDD.t0 DVDD.t367 56.231
R2484 DVDD.t202 DVDD.t292 56.231
R2485 DVDD.t494 DVDD.t394 56.231
R2486 DVDD.t329 DVDD.t411 56.231
R2487 DVDD.t182 DVDD.t184 56.231
R2488 DVDD.t465 DVDD.t108 56.231
R2489 DVDD.t217 DVDD.t408 56.231
R2490 DVDD.t50 DVDD.t488 56.231
R2491 DVDD.t168 DVDD.t472 56.231
R2492 DVDD.t233 DVDD.t391 56.231
R2493 DVDD.t365 DVDD.t115 56.231
R2494 DVDD.t102 DVDD.t188 56.231
R2495 DVDD.t210 DVDD.t386 56.231
R2496 DVDD.t272 DVDD.t306 56.231
R2497 DVDD.t515 DVDD.t27 56.231
R2498 DVDD.t502 DVDD.t166 56.231
R2499 DVDD.t187 DVDD.t134 54.7513
R2500 DVDD.t393 DVDD.t399 54.7513
R2501 DVDD.t197 DVDD.t506 54.7513
R2502 DVDD.t526 DVDD.t37 54.7513
R2503 DVDD.t238 DVDD.t252 45.8728
R2504 DVDD.t350 DVDD.t124 45.8728
R2505 DVDD.t396 DVDD.t132 45.8728
R2506 DVDD.t259 DVDD.t111 45.8728
R2507 DVDD.t215 DVDD.t20 45.8728
R2508 DVDD.t485 DVDD.t321 45.8728
R2509 DVDD.n745 DVDD.n744 43.9358
R2510 DVDD.n779 DVDD.n778 43.9358
R2511 DVDD.n128 DVDD.n127 43.9358
R2512 DVDD.n769 DVDD.n144 43.9358
R2513 DVDD.n101 DVDD.n98 43.9358
R2514 DVDD.n813 DVDD.n812 43.9358
R2515 DVDD.n91 DVDD.n90 43.9358
R2516 DVDD.n702 DVDD.n486 43.9358
R2517 DVDD.n669 DVDD.n668 43.9358
R2518 DVDD.n544 DVDD.n517 43.9358
R2519 DVDD.n602 DVDD.n569 43.9358
R2520 DVDD.n659 DVDD.n641 43.9358
R2521 DVDD.n678 DVDD.n677 43.9358
R2522 DVDD.n535 DVDD.n521 43.9358
R2523 DVDD.n553 DVDD.n552 43.9358
R2524 DVDD.n453 DVDD.n179 43.9358
R2525 DVDD.n422 DVDD.n421 43.9358
R2526 DVDD.n412 DVDD.n394 43.9358
R2527 DVDD.n228 DVDD.n202 43.9358
R2528 DVDD.n366 DVDD.n253 43.9358
R2529 DVDD.n237 DVDD.n236 43.9358
R2530 DVDD.n622 DVDD.n497 43.1829
R2531 DVDD.n621 DVDD.n620 43.1829
R2532 DVDD.n305 DVDD.n304 43.1829
R2533 DVDD.n303 DVDD.n302 43.1829
R2534 DVDD.n733 DVDD.n167 42.302
R2535 DVDD.n760 DVDD.n759 42.302
R2536 DVDD.n80 DVDD.n78 42.302
R2537 DVDD.n827 DVDD.n37 42.302
R2538 DVDD.n720 DVDD.n478 42.302
R2539 DVDD.n650 DVDD.n649 42.302
R2540 DVDD.n566 DVDD.n504 42.302
R2541 DVDD.n585 DVDD.n584 42.302
R2542 DVDD.n471 DVDD.n171 42.302
R2543 DVDD.n403 DVDD.n402 42.302
R2544 DVDD.n250 DVDD.n189 42.302
R2545 DVDD.n349 DVDD.n348 42.302
R2546 DVDD.n166 DVDD.n162 41.549
R2547 DVDD.n821 DVDD.n820 41.549
R2548 DVDD.n709 DVDD.n482 41.549
R2549 DVDD.n595 DVDD.n575 41.549
R2550 DVDD.n460 DVDD.n175 41.549
R2551 DVDD.n359 DVDD.n259 41.549
R2552 DVDD.n330 DVDD.n324 41.5414
R2553 DVDD.n318 DVDD.n317 41.5414
R2554 DVDD.n290 DVDD.n284 41.5414
R2555 DVDD.n338 DVDD.n337 41.5414
R2556 DVDD.t336 DVDD.t304 36.9943
R2557 DVDD.t40 DVDD.t249 36.9943
R2558 DVDD.n691 DVDD.t356 36.9943
R2559 DVDD.n614 DVDD.t446 36.9943
R2560 DVDD.t89 DVDD.t455 36.9943
R2561 DVDD.t223 DVDD.t285 36.9943
R2562 DVDD.n328 DVDD.n327 34.6358
R2563 DVDD.n789 DVDD.n135 34.6358
R2564 DVDD.n736 DVDD.n735 34.6358
R2565 DVDD.n767 DVDD.n147 34.6358
R2566 DVDD.n112 DVDD.n111 34.6358
R2567 DVDD.n88 DVDD.n71 34.6358
R2568 DVDD.n823 DVDD.n822 34.6358
R2569 DVDD.n168 DVDD.n163 34.6358
R2570 DVDD.n169 DVDD.n168 34.6358
R2571 DVDD.n730 DVDD.n169 34.6358
R2572 DVDD.n740 DVDD.n739 34.6358
R2573 DVDD.n756 DVDD.n153 34.6358
R2574 DVDD.n749 DVDD.n153 34.6358
R2575 DVDD.n749 DVDD.n748 34.6358
R2576 DVDD.n772 DVDD.n143 34.6358
R2577 DVDD.n764 DVDD.n143 34.6358
R2578 DVDD.n764 DVDD.n763 34.6358
R2579 DVDD.n776 DVDD.n775 34.6358
R2580 DVDD.n792 DVDD.n133 34.6358
R2581 DVDD.n785 DVDD.n133 34.6358
R2582 DVDD.n785 DVDD.n784 34.6358
R2583 DVDD.n107 DVDD.n106 34.6358
R2584 DVDD.n107 DVDD.n60 34.6358
R2585 DVDD.n115 DVDD.n60 34.6358
R2586 DVDD.n96 DVDD.n95 34.6358
R2587 DVDD.n84 DVDD.n83 34.6358
R2588 DVDD.n84 DVDD.n68 34.6358
R2589 DVDD.n93 DVDD.n68 34.6358
R2590 DVDD.n809 DVDD.n808 34.6358
R2591 DVDD.n808 DVDD.n53 34.6358
R2592 DVDD.n75 DVDD.n53 34.6358
R2593 DVDD.n818 DVDD.n817 34.6358
R2594 DVDD.n39 DVDD.n38 34.6358
R2595 DVDD.n40 DVDD.n39 34.6358
R2596 DVDD.n46 DVDD.n40 34.6358
R2597 DVDD.n718 DVDD.n717 34.6358
R2598 DVDD.n657 DVDD.n644 34.6358
R2599 DVDD.n625 DVDD.n624 34.6358
R2600 DVDD.n687 DVDD.n625 34.6358
R2601 DVDD.n687 DVDD.n686 34.6358
R2602 DVDD.n686 DVDD.n685 34.6358
R2603 DVDD.n685 DVDD.n626 34.6358
R2604 DVDD.n533 DVDD.n524 34.6358
R2605 DVDD.n527 DVDD.n524 34.6358
R2606 DVDD.n527 DVDD.n500 34.6358
R2607 DVDD.n618 DVDD.n500 34.6358
R2608 DVDD.n619 DVDD.n618 34.6358
R2609 DVDD.n560 DVDD.n559 34.6358
R2610 DVDD.n588 DVDD.n587 34.6358
R2611 DVDD.n715 DVDD.n714 34.6358
R2612 DVDD.n714 DVDD.n479 34.6358
R2613 DVDD.n723 DVDD.n479 34.6358
R2614 DVDD.n712 DVDD.n711 34.6358
R2615 DVDD.n697 DVDD.n696 34.6358
R2616 DVDD.n697 DVDD.n489 34.6358
R2617 DVDD.n705 DVDD.n489 34.6358
R2618 DVDD.n662 DVDD.n640 34.6358
R2619 DVDD.n654 DVDD.n640 34.6358
R2620 DVDD.n654 DVDD.n653 34.6358
R2621 DVDD.n666 DVDD.n665 34.6358
R2622 DVDD.n681 DVDD.n629 34.6358
R2623 DVDD.n675 DVDD.n629 34.6358
R2624 DVDD.n675 DVDD.n674 34.6358
R2625 DVDD.n540 DVDD.n539 34.6358
R2626 DVDD.n539 DVDD.n538 34.6358
R2627 DVDD.n538 DVDD.n520 34.6358
R2628 DVDD.n550 DVDD.n549 34.6358
R2629 DVDD.n563 DVDD.n506 34.6358
R2630 DVDD.n556 DVDD.n506 34.6358
R2631 DVDD.n556 DVDD.n555 34.6358
R2632 DVDD.n570 DVDD.n567 34.6358
R2633 DVDD.n607 DVDD.n567 34.6358
R2634 DVDD.n608 DVDD.n607 34.6358
R2635 DVDD.n593 DVDD.n573 34.6358
R2636 DVDD.n582 DVDD.n578 34.6358
R2637 DVDD.n590 DVDD.n578 34.6358
R2638 DVDD.n591 DVDD.n590 34.6358
R2639 DVDD.n432 DVDD.n385 34.6358
R2640 DVDD.n469 DVDD.n468 34.6358
R2641 DVDD.n410 DVDD.n397 34.6358
R2642 DVDD.n219 DVDD.n218 34.6358
R2643 DVDD.n244 DVDD.n243 34.6358
R2644 DVDD.n352 DVDD.n351 34.6358
R2645 DVDD.n466 DVDD.n465 34.6358
R2646 DVDD.n465 DVDD.n172 34.6358
R2647 DVDD.n474 DVDD.n172 34.6358
R2648 DVDD.n463 DVDD.n462 34.6358
R2649 DVDD.n448 DVDD.n447 34.6358
R2650 DVDD.n448 DVDD.n182 34.6358
R2651 DVDD.n456 DVDD.n182 34.6358
R2652 DVDD.n415 DVDD.n393 34.6358
R2653 DVDD.n407 DVDD.n393 34.6358
R2654 DVDD.n407 DVDD.n406 34.6358
R2655 DVDD.n419 DVDD.n418 34.6358
R2656 DVDD.n435 DVDD.n383 34.6358
R2657 DVDD.n428 DVDD.n383 34.6358
R2658 DVDD.n428 DVDD.n427 34.6358
R2659 DVDD.n224 DVDD.n223 34.6358
R2660 DVDD.n223 DVDD.n222 34.6358
R2661 DVDD.n222 DVDD.n205 34.6358
R2662 DVDD.n234 DVDD.n233 34.6358
R2663 DVDD.n247 DVDD.n191 34.6358
R2664 DVDD.n240 DVDD.n191 34.6358
R2665 DVDD.n240 DVDD.n239 34.6358
R2666 DVDD.n254 DVDD.n251 34.6358
R2667 DVDD.n371 DVDD.n251 34.6358
R2668 DVDD.n372 DVDD.n371 34.6358
R2669 DVDD.n357 DVDD.n257 34.6358
R2670 DVDD.n346 DVDD.n262 34.6358
R2671 DVDD.n354 DVDD.n262 34.6358
R2672 DVDD.n355 DVDD.n354 34.6358
R2673 DVDD.n320 DVDD.n319 34.6358
R2674 DVDD.n307 DVDD.n306 34.6358
R2675 DVDD.n307 DVDD.n274 34.6358
R2676 DVDD.n311 DVDD.n274 34.6358
R2677 DVDD.n312 DVDD.n311 34.6358
R2678 DVDD.n313 DVDD.n312 34.6358
R2679 DVDD.n295 DVDD.n294 34.6358
R2680 DVDD.n296 DVDD.n295 34.6358
R2681 DVDD.n296 DVDD.n279 34.6358
R2682 DVDD.n300 DVDD.n279 34.6358
R2683 DVDD.n301 DVDD.n300 34.6358
R2684 DVDD.n288 DVDD.n287 34.6358
R2685 DVDD.n340 DVDD.n339 34.6358
R2686 DVDD.n920 DVDD.n2 34.6358
R2687 DVDD.n921 DVDD.n920 34.6358
R2688 DVDD.n923 DVDD.n921 34.6358
R2689 DVDD.n916 DVDD.n913 34.6358
R2690 DVDD.n905 DVDD.n7 34.6358
R2691 DVDD.n906 DVDD.n905 34.6358
R2692 DVDD.n907 DVDD.n906 34.6358
R2693 DVDD.n893 DVDD.n9 34.6358
R2694 DVDD.n897 DVDD.n9 34.6358
R2695 DVDD.n898 DVDD.n897 34.6358
R2696 DVDD.n891 DVDD.n890 34.6358
R2697 DVDD.n881 DVDD.n880 34.6358
R2698 DVDD.n881 DVDD.n15 34.6358
R2699 DVDD.n885 DVDD.n15 34.6358
R2700 DVDD.n868 DVDD.n18 34.6358
R2701 DVDD.n872 DVDD.n18 34.6358
R2702 DVDD.n873 DVDD.n872 34.6358
R2703 DVDD.n863 DVDD.n862 34.6358
R2704 DVDD.n856 DVDD.n855 34.6358
R2705 DVDD.n856 DVDD.n24 34.6358
R2706 DVDD.n860 DVDD.n24 34.6358
R2707 DVDD.n845 DVDD.n27 34.6358
R2708 DVDD.n849 DVDD.n27 34.6358
R2709 DVDD.n850 DVDD.n849 34.6358
R2710 DVDD.n840 DVDD.n839 34.6358
R2711 DVDD.n833 DVDD.n832 34.6358
R2712 DVDD.n833 DVDD.n33 34.6358
R2713 DVDD.n837 DVDD.n33 34.6358
R2714 DVDD.n769 DVDD.n768 33.8829
R2715 DVDD.n90 DVDD.n89 33.8829
R2716 DVDD.n659 DVDD.n658 33.8829
R2717 DVDD.n552 DVDD.n510 33.8829
R2718 DVDD.n412 DVDD.n411 33.8829
R2719 DVDD.n236 DVDD.n195 33.8829
R2720 DVDD.n742 DVDD.n156 32.7534
R2721 DVDD.n783 DVDD.n137 32.7534
R2722 DVDD.n105 DVDD.n104 32.7534
R2723 DVDD.n815 DVDD.n49 32.7534
R2724 DVDD.n707 DVDD.n706 32.7534
R2725 DVDD.n673 DVDD.n634 32.7534
R2726 DVDD.n547 DVDD.n516 32.7534
R2727 DVDD.n599 DVDD.n598 32.7534
R2728 DVDD.n458 DVDD.n457 32.7534
R2729 DVDD.n426 DVDD.n387 32.7534
R2730 DVDD.n231 DVDD.n201 32.7534
R2731 DVDD.n363 DVDD.n362 32.7534
R2732 DVDD.n911 DVDD.n5 32.7534
R2733 DVDD.n887 DVDD.n886 32.7534
R2734 DVDD.n867 DVDD.n866 32.7534
R2735 DVDD.n844 DVDD.n843 32.7534
R2736 DVDD.t352 DVDD.t54 31.0753
R2737 DVDD.t354 DVDD.t296 31.0753
R2738 DVDD.t328 DVDD.t448 31.0753
R2739 DVDD.t359 DVDD.t510 31.0753
R2740 DVDD.n796 DVDD.n131 30.8711
R2741 DVDD.n119 DVDD.n58 30.8711
R2742 DVDD.n439 DVDD.n381 30.8711
R2743 DVDD.n212 DVDD.n210 30.8711
R2744 DVDD.n757 DVDD.n756 29.7417
R2745 DVDD.n793 DVDD.n792 29.7417
R2746 DVDD.n116 DVDD.n115 29.7417
R2747 DVDD.n76 DVDD.n75 29.7417
R2748 DVDD.n696 DVDD.n491 29.7417
R2749 DVDD.n682 DVDD.n681 29.7417
R2750 DVDD.n530 DVDD.n520 29.7417
R2751 DVDD.n609 DVDD.n608 29.7417
R2752 DVDD.n447 DVDD.n184 29.7417
R2753 DVDD.n436 DVDD.n435 29.7417
R2754 DVDD.n215 DVDD.n205 29.7417
R2755 DVDD.n373 DVDD.n372 29.7417
R2756 DVDD.n901 DVDD.n7 29.7417
R2757 DVDD.n880 DVDD.n879 29.7417
R2758 DVDD.n874 DVDD.n873 29.7417
R2759 DVDD.n851 DVDD.n850 29.7417
R2760 DVDD.n496 DVDD.t120 28.752
R2761 DVDD.n499 DVDD.t378 28.752
R2762 DVDD.n276 DVDD.t52 28.752
R2763 DVDD.n278 DVDD.t327 28.752
R2764 DVDD.n327 DVDD.n326 27.8593
R2765 DVDD.n735 DVDD.n734 27.8593
R2766 DVDD.n151 DVDD.n147 27.8593
R2767 DVDD.n79 DVDD.n71 27.8593
R2768 DVDD.n823 DVDD.n42 27.8593
R2769 DVDD.n719 DVDD.n718 27.8593
R2770 DVDD.n648 DVDD.n644 27.8593
R2771 DVDD.n560 DVDD.n508 27.8593
R2772 DVDD.n588 DVDD.n586 27.8593
R2773 DVDD.n470 DVDD.n469 27.8593
R2774 DVDD.n401 DVDD.n397 27.8593
R2775 DVDD.n244 DVDD.n193 27.8593
R2776 DVDD.n352 DVDD.n350 27.8593
R2777 DVDD.n320 DVDD.n268 27.8593
R2778 DVDD.n287 DVDD.n286 27.8593
R2779 DVDD.n340 DVDD.n264 27.8593
R2780 DVDD.n753 DVDD.n152 26.6181
R2781 DVDD.n754 DVDD.n753 26.6181
R2782 DVDD.n800 DVDD.n123 26.6181
R2783 DVDD.n800 DVDD.n799 26.6181
R2784 DVDD.n805 DVDD.n804 26.6181
R2785 DVDD.n804 DVDD.n55 26.6181
R2786 DVDD.n612 DVDD.n502 26.6181
R2787 DVDD.n612 DVDD.n611 26.6181
R2788 DVDD.n694 DVDD.n693 26.6181
R2789 DVDD.n693 DVDD.n490 26.6181
R2790 DVDD.n690 DVDD.n493 26.6181
R2791 DVDD.n690 DVDD.n689 26.6181
R2792 DVDD.n615 DVDD.n501 26.6181
R2793 DVDD.n616 DVDD.n615 26.6181
R2794 DVDD.n445 DVDD.n444 26.6181
R2795 DVDD.n444 DVDD.n183 26.6181
R2796 DVDD.n376 DVDD.n187 26.6181
R2797 DVDD.n376 DVDD.n375 26.6181
R2798 DVDD.n323 DVDD.t122 26.5955
R2799 DVDD.n323 DVDD.t101 26.5955
R2800 DVDD.n130 DVDD.t305 26.5955
R2801 DVDD.n130 DVDD.t135 26.5955
R2802 DVDD.n165 DVDD.t97 26.5955
R2803 DVDD.n165 DVDD.t288 26.5955
R2804 DVDD.n146 DVDD.t418 26.5955
R2805 DVDD.n146 DVDD.t425 26.5955
R2806 DVDD.n57 DVDD.t400 26.5955
R2807 DVDD.n57 DVDD.t250 26.5955
R2808 DVDD.n70 DVDD.t84 26.5955
R2809 DVDD.n70 DVDD.t154 26.5955
R2810 DVDD.n43 DVDD.t395 26.5955
R2811 DVDD.n43 DVDD.t412 26.5955
R2812 DVDD.n481 DVDD.t185 26.5955
R2813 DVDD.n481 DVDD.t109 26.5955
R2814 DVDD.n643 DVDD.t86 26.5955
R2815 DVDD.n643 DVDD.t105 26.5955
R2816 DVDD.n509 DVDD.t341 26.5955
R2817 DVDD.n509 DVDD.t227 26.5955
R2818 DVDD.n574 DVDD.t473 26.5955
R2819 DVDD.n574 DVDD.t392 26.5955
R2820 DVDD.n380 DVDD.t456 26.5955
R2821 DVDD.n380 DVDD.t507 26.5955
R2822 DVDD.n174 DVDD.t116 26.5955
R2823 DVDD.n174 DVDD.t189 26.5955
R2824 DVDD.n396 DVDD.t372 26.5955
R2825 DVDD.n396 DVDD.t32 26.5955
R2826 DVDD.n209 DVDD.t527 26.5955
R2827 DVDD.n209 DVDD.t224 26.5955
R2828 DVDD.n194 DVDD.t173 26.5955
R2829 DVDD.n194 DVDD.t343 26.5955
R2830 DVDD.n258 DVDD.t28 26.5955
R2831 DVDD.n258 DVDD.t167 26.5955
R2832 DVDD.n270 DVDD.t88 26.5955
R2833 DVDD.n270 DVDD.t92 26.5955
R2834 DVDD.n283 DVDD.t282 26.5955
R2835 DVDD.n283 DVDD.t280 26.5955
R2836 DVDD.n266 DVDD.t45 26.5955
R2837 DVDD.n266 DVDD.t274 26.5955
R2838 DVDD.n797 DVDD.n796 25.977
R2839 DVDD.n120 DVDD.n119 25.977
R2840 DVDD.n440 DVDD.n439 25.977
R2841 DVDD.n212 DVDD.n211 25.977
R2842 DVDD.n315 DVDD.n272 24.9767
R2843 DVDD.n292 DVDD.n282 24.9767
R2844 DVDD.n793 DVDD.n129 23.9829
R2845 DVDD.n116 DVDD.n56 23.9829
R2846 DVDD.n682 DVDD.n627 23.9829
R2847 DVDD.n530 DVDD.n529 23.9829
R2848 DVDD.n436 DVDD.n379 23.9829
R2849 DVDD.n215 DVDD.n214 23.9829
R2850 DVDD.n789 DVDD.n788 22.9652
R2851 DVDD.n112 DVDD.n110 22.9652
R2852 DVDD.n432 DVDD.n431 22.9652
R2853 DVDD.n219 DVDD.n208 22.9652
R2854 DVDD.t251 DVDD.t319 19.2373
R2855 DVDD.t127 DVDD.t450 19.2373
R2856 DVDD.t22 DVDD.t468 19.2373
R2857 DVDD.t198 DVDD.t484 19.2373
R2858 DVDD.t73 DVDD.t361 17.7575
R2859 DVDD.t228 DVDD.t517 17.7575
R2860 DVDD.t206 DVDD.t204 17.7575
R2861 DVDD.t76 DVDD.t402 17.7575
R2862 DVDD.t388 DVDD.t384 17.7575
R2863 DVDD.t522 DVDD.t277 17.7575
R2864 DVDD.n158 DVDD.n154 17.5829
R2865 DVDD.n140 DVDD.n138 17.5829
R2866 DVDD.n125 DVDD.n124 17.5829
R2867 DVDD.n100 DVDD.n99 17.5829
R2868 DVDD.n52 DVDD.n51 17.5829
R2869 DVDD.n701 DVDD.n700 17.5829
R2870 DVDD.n637 DVDD.n635 17.5829
R2871 DVDD.n543 DVDD.n542 17.5829
R2872 DVDD.n604 DVDD.n603 17.5829
R2873 DVDD.n452 DVDD.n451 17.5829
R2874 DVDD.n390 DVDD.n388 17.5829
R2875 DVDD.n227 DVDD.n226 17.5829
R2876 DVDD.n368 DVDD.n367 17.5829
R2877 DVDD.n632 DVDD.n626 17.3181
R2878 DVDD.n678 DVDD.n632 17.3181
R2879 DVDD.n535 DVDD.n534 17.3181
R2880 DVDD.n534 DVDD.n533 17.3181
R2881 DVDD.n313 DVDD.n272 17.3181
R2882 DVDD.n294 DVDD.n282 17.3181
R2883 DVDD.n729 DVDD.n728 16.077
R2884 DVDD.n150 DVDD.n149 16.077
R2885 DVDD.n74 DVDD.n73 16.077
R2886 DVDD.n828 DVDD.n36 16.077
R2887 DVDD.n725 DVDD.n724 16.077
R2888 DVDD.n647 DVDD.n646 16.077
R2889 DVDD.n565 DVDD.n564 16.077
R2890 DVDD.n581 DVDD.n580 16.077
R2891 DVDD.n476 DVDD.n475 16.077
R2892 DVDD.n400 DVDD.n399 16.077
R2893 DVDD.n249 DVDD.n248 16.077
R2894 DVDD.n345 DVDD.n344 16.077
R2895 DVDD.n922 DVDD.n1 16.077
R2896 DVDD.n900 DVDD.n899 16.077
R2897 DVDD.n854 DVDD.n853 16.077
R2898 DVDD.n831 DVDD.n830 16.077
R2899 DVDD.n326 DVDD.n170 14.3803
R2900 DVDD.n322 DVDD.n268 14.3803
R2901 DVDD.n286 DVDD.n267 14.3803
R2902 DVDD.n342 DVDD.n264 14.3803
R2903 DVDD.t78 DVDD.t106 13.3183
R2904 DVDD.t347 DVDD.t492 13.3183
R2905 DVDD.t373 DVDD.t499 13.3183
R2906 DVDD.t529 DVDD.t10 13.3183
R2907 DVDD.t314 DVDD.t61 13.3183
R2908 DVDD.t195 DVDD.t140 13.3183
R2909 DVDD.n748 DVDD.n156 11.6711
R2910 DVDD.n784 DVDD.n783 11.6711
R2911 DVDD.n106 DVDD.n105 11.6711
R2912 DVDD.n809 DVDD.n49 11.6711
R2913 DVDD.n706 DVDD.n705 11.6711
R2914 DVDD.n674 DVDD.n673 11.6711
R2915 DVDD.n540 DVDD.n516 11.6711
R2916 DVDD.n599 DVDD.n570 11.6711
R2917 DVDD.n457 DVDD.n456 11.6711
R2918 DVDD.n427 DVDD.n426 11.6711
R2919 DVDD.n224 DVDD.n201 11.6711
R2920 DVDD.n363 DVDD.n254 11.6711
R2921 DVDD.n907 DVDD.n5 11.6711
R2922 DVDD.n886 DVDD.n885 11.6711
R2923 DVDD.n868 DVDD.n867 11.6711
R2924 DVDD.n845 DVDD.n844 11.6711
R2925 DVDD.n745 DVDD.n158 10.5417
R2926 DVDD.n779 DVDD.n140 10.5417
R2927 DVDD.n127 DVDD.n124 10.5417
R2928 DVDD.n101 DVDD.n100 10.5417
R2929 DVDD.n812 DVDD.n51 10.5417
R2930 DVDD.n702 DVDD.n701 10.5417
R2931 DVDD.n669 DVDD.n637 10.5417
R2932 DVDD.n544 DVDD.n543 10.5417
R2933 DVDD.n603 DVDD.n602 10.5417
R2934 DVDD.n453 DVDD.n452 10.5417
R2935 DVDD.n422 DVDD.n390 10.5417
R2936 DVDD.n228 DVDD.n227 10.5417
R2937 DVDD.n367 DVDD.n366 10.5417
R2938 DVDD.n826 DVDD.n38 9.3005
R2939 DVDD.n825 DVDD.n39 9.3005
R2940 DVDD.n824 DVDD.n40 9.3005
R2941 DVDD.n46 DVDD.n41 9.3005
R2942 DVDD.n819 DVDD.n818 9.3005
R2943 DVDD.n817 DVDD.n44 9.3005
R2944 DVDD.n815 DVDD.n814 9.3005
R2945 DVDD.n50 DVDD.n49 9.3005
R2946 DVDD.n810 DVDD.n809 9.3005
R2947 DVDD.n808 DVDD.n807 9.3005
R2948 DVDD.n806 DVDD.n53 9.3005
R2949 DVDD.n75 DVDD.n54 9.3005
R2950 DVDD.n83 DVDD.n82 9.3005
R2951 DVDD.n85 DVDD.n84 9.3005
R2952 DVDD.n86 DVDD.n68 9.3005
R2953 DVDD.n93 DVDD.n92 9.3005
R2954 DVDD.n95 DVDD.n66 9.3005
R2955 DVDD.n97 DVDD.n96 9.3005
R2956 DVDD.n104 DVDD.n103 9.3005
R2957 DVDD.n105 DVDD.n63 9.3005
R2958 DVDD.n106 DVDD.n62 9.3005
R2959 DVDD.n108 DVDD.n107 9.3005
R2960 DVDD.n61 DVDD.n60 9.3005
R2961 DVDD.n115 DVDD.n114 9.3005
R2962 DVDD.n117 DVDD.n116 9.3005
R2963 DVDD.n794 DVDD.n793 9.3005
R2964 DVDD.n792 DVDD.n791 9.3005
R2965 DVDD.n134 DVDD.n133 9.3005
R2966 DVDD.n786 DVDD.n785 9.3005
R2967 DVDD.n784 DVDD.n136 9.3005
R2968 DVDD.n783 DVDD.n781 9.3005
R2969 DVDD.n139 DVDD.n137 9.3005
R2970 DVDD.n777 DVDD.n776 9.3005
R2971 DVDD.n775 DVDD.n141 9.3005
R2972 DVDD.n772 DVDD.n771 9.3005
R2973 DVDD.n145 DVDD.n143 9.3005
R2974 DVDD.n765 DVDD.n764 9.3005
R2975 DVDD.n763 DVDD.n762 9.3005
R2976 DVDD.n756 DVDD.n755 9.3005
R2977 DVDD.n751 DVDD.n153 9.3005
R2978 DVDD.n750 DVDD.n749 9.3005
R2979 DVDD.n748 DVDD.n747 9.3005
R2980 DVDD.n157 DVDD.n156 9.3005
R2981 DVDD.n743 DVDD.n742 9.3005
R2982 DVDD.n740 DVDD.n159 9.3005
R2983 DVDD.n739 DVDD.n738 9.3005
R2984 DVDD.n737 DVDD.n163 9.3005
R2985 DVDD.n168 DVDD.n164 9.3005
R2986 DVDD.n732 DVDD.n169 9.3005
R2987 DVDD.n731 DVDD.n730 9.3005
R2988 DVDD.n825 DVDD.n37 9.3005
R2989 DVDD.n824 DVDD.n823 9.3005
R2990 DVDD.n822 DVDD.n41 9.3005
R2991 DVDD.n90 DVDD.n69 9.3005
R2992 DVDD.n81 DVDD.n80 9.3005
R2993 DVDD.n72 DVDD.n71 9.3005
R2994 DVDD.n88 DVDD.n87 9.3005
R2995 DVDD.n812 DVDD.n811 9.3005
R2996 DVDD.n102 DVDD.n101 9.3005
R2997 DVDD.n121 DVDD.n120 9.3005
R2998 DVDD.n110 DVDD.n109 9.3005
R2999 DVDD.n113 DVDD.n112 9.3005
R3000 DVDD.n111 DVDD.n59 9.3005
R3001 DVDD.n119 DVDD.n118 9.3005
R3002 DVDD.n761 DVDD.n760 9.3005
R3003 DVDD.n770 DVDD.n769 9.3005
R3004 DVDD.n767 DVDD.n766 9.3005
R3005 DVDD.n148 DVDD.n147 9.3005
R3006 DVDD.n733 DVDD.n732 9.3005
R3007 DVDD.n737 DVDD.n736 9.3005
R3008 DVDD.n735 DVDD.n164 9.3005
R3009 DVDD.n127 DVDD.n126 9.3005
R3010 DVDD.n788 DVDD.n787 9.3005
R3011 DVDD.n790 DVDD.n789 9.3005
R3012 DVDD.n135 DVDD.n132 9.3005
R3013 DVDD.n796 DVDD.n795 9.3005
R3014 DVDD.n798 DVDD.n797 9.3005
R3015 DVDD.n780 DVDD.n779 9.3005
R3016 DVDD.n746 DVDD.n745 9.3005
R3017 DVDD.n583 DVDD.n582 9.3005
R3018 DVDD.n579 DVDD.n578 9.3005
R3019 DVDD.n590 DVDD.n589 9.3005
R3020 DVDD.n591 DVDD.n576 9.3005
R3021 DVDD.n594 DVDD.n593 9.3005
R3022 DVDD.n596 DVDD.n573 9.3005
R3023 DVDD.n598 DVDD.n597 9.3005
R3024 DVDD.n600 DVDD.n599 9.3005
R3025 DVDD.n570 DVDD.n568 9.3005
R3026 DVDD.n605 DVDD.n567 9.3005
R3027 DVDD.n607 DVDD.n606 9.3005
R3028 DVDD.n608 DVDD.n503 9.3005
R3029 DVDD.n563 DVDD.n562 9.3005
R3030 DVDD.n507 DVDD.n506 9.3005
R3031 DVDD.n557 DVDD.n556 9.3005
R3032 DVDD.n555 DVDD.n554 9.3005
R3033 DVDD.n551 DVDD.n550 9.3005
R3034 DVDD.n549 DVDD.n514 9.3005
R3035 DVDD.n547 DVDD.n546 9.3005
R3036 DVDD.n518 DVDD.n516 9.3005
R3037 DVDD.n541 DVDD.n540 9.3005
R3038 DVDD.n539 DVDD.n519 9.3005
R3039 DVDD.n538 DVDD.n537 9.3005
R3040 DVDD.n522 DVDD.n520 9.3005
R3041 DVDD.n531 DVDD.n530 9.3005
R3042 DVDD.n683 DVDD.n682 9.3005
R3043 DVDD.n681 DVDD.n680 9.3005
R3044 DVDD.n630 DVDD.n629 9.3005
R3045 DVDD.n676 DVDD.n675 9.3005
R3046 DVDD.n674 DVDD.n633 9.3005
R3047 DVDD.n673 DVDD.n671 9.3005
R3048 DVDD.n636 DVDD.n634 9.3005
R3049 DVDD.n667 DVDD.n666 9.3005
R3050 DVDD.n665 DVDD.n638 9.3005
R3051 DVDD.n662 DVDD.n661 9.3005
R3052 DVDD.n642 DVDD.n640 9.3005
R3053 DVDD.n655 DVDD.n654 9.3005
R3054 DVDD.n653 DVDD.n652 9.3005
R3055 DVDD.n696 DVDD.n695 9.3005
R3056 DVDD.n698 DVDD.n697 9.3005
R3057 DVDD.n699 DVDD.n489 9.3005
R3058 DVDD.n705 DVDD.n704 9.3005
R3059 DVDD.n706 DVDD.n487 9.3005
R3060 DVDD.n708 DVDD.n707 9.3005
R3061 DVDD.n711 DVDD.n710 9.3005
R3062 DVDD.n712 DVDD.n483 9.3005
R3063 DVDD.n716 DVDD.n715 9.3005
R3064 DVDD.n714 DVDD.n480 9.3005
R3065 DVDD.n721 DVDD.n479 9.3005
R3066 DVDD.n723 DVDD.n722 9.3005
R3067 DVDD.n585 DVDD.n579 9.3005
R3068 DVDD.n589 DVDD.n588 9.3005
R3069 DVDD.n587 DVDD.n576 9.3005
R3070 DVDD.n552 DVDD.n511 9.3005
R3071 DVDD.n505 DVDD.n504 9.3005
R3072 DVDD.n561 DVDD.n560 9.3005
R3073 DVDD.n559 DVDD.n558 9.3005
R3074 DVDD.n536 DVDD.n535 9.3005
R3075 DVDD.n533 DVDD.n532 9.3005
R3076 DVDD.n525 DVDD.n524 9.3005
R3077 DVDD.n528 DVDD.n527 9.3005
R3078 DVDD.n526 DVDD.n500 9.3005
R3079 DVDD.n618 DVDD.n617 9.3005
R3080 DVDD.n619 DVDD.n498 9.3005
R3081 DVDD.n679 DVDD.n678 9.3005
R3082 DVDD.n624 DVDD.n623 9.3005
R3083 DVDD.n625 DVDD.n494 9.3005
R3084 DVDD.n688 DVDD.n687 9.3005
R3085 DVDD.n686 DVDD.n495 9.3005
R3086 DVDD.n685 DVDD.n684 9.3005
R3087 DVDD.n628 DVDD.n626 9.3005
R3088 DVDD.n651 DVDD.n650 9.3005
R3089 DVDD.n660 DVDD.n659 9.3005
R3090 DVDD.n657 DVDD.n656 9.3005
R3091 DVDD.n645 DVDD.n644 9.3005
R3092 DVDD.n721 DVDD.n720 9.3005
R3093 DVDD.n717 DVDD.n716 9.3005
R3094 DVDD.n718 DVDD.n480 9.3005
R3095 DVDD.n602 DVDD.n601 9.3005
R3096 DVDD.n545 DVDD.n544 9.3005
R3097 DVDD.n670 DVDD.n669 9.3005
R3098 DVDD.n703 DVDD.n702 9.3005
R3099 DVDD.n347 DVDD.n346 9.3005
R3100 DVDD.n263 DVDD.n262 9.3005
R3101 DVDD.n354 DVDD.n353 9.3005
R3102 DVDD.n355 DVDD.n260 9.3005
R3103 DVDD.n358 DVDD.n357 9.3005
R3104 DVDD.n360 DVDD.n257 9.3005
R3105 DVDD.n362 DVDD.n361 9.3005
R3106 DVDD.n364 DVDD.n363 9.3005
R3107 DVDD.n254 DVDD.n252 9.3005
R3108 DVDD.n369 DVDD.n251 9.3005
R3109 DVDD.n371 DVDD.n370 9.3005
R3110 DVDD.n372 DVDD.n188 9.3005
R3111 DVDD.n247 DVDD.n246 9.3005
R3112 DVDD.n192 DVDD.n191 9.3005
R3113 DVDD.n241 DVDD.n240 9.3005
R3114 DVDD.n239 DVDD.n238 9.3005
R3115 DVDD.n235 DVDD.n234 9.3005
R3116 DVDD.n233 DVDD.n199 9.3005
R3117 DVDD.n231 DVDD.n230 9.3005
R3118 DVDD.n203 DVDD.n201 9.3005
R3119 DVDD.n225 DVDD.n224 9.3005
R3120 DVDD.n223 DVDD.n204 9.3005
R3121 DVDD.n222 DVDD.n221 9.3005
R3122 DVDD.n207 DVDD.n205 9.3005
R3123 DVDD.n216 DVDD.n215 9.3005
R3124 DVDD.n437 DVDD.n436 9.3005
R3125 DVDD.n435 DVDD.n434 9.3005
R3126 DVDD.n384 DVDD.n383 9.3005
R3127 DVDD.n429 DVDD.n428 9.3005
R3128 DVDD.n427 DVDD.n386 9.3005
R3129 DVDD.n426 DVDD.n424 9.3005
R3130 DVDD.n389 DVDD.n387 9.3005
R3131 DVDD.n420 DVDD.n419 9.3005
R3132 DVDD.n418 DVDD.n391 9.3005
R3133 DVDD.n415 DVDD.n414 9.3005
R3134 DVDD.n395 DVDD.n393 9.3005
R3135 DVDD.n408 DVDD.n407 9.3005
R3136 DVDD.n406 DVDD.n405 9.3005
R3137 DVDD.n447 DVDD.n446 9.3005
R3138 DVDD.n449 DVDD.n448 9.3005
R3139 DVDD.n450 DVDD.n182 9.3005
R3140 DVDD.n456 DVDD.n455 9.3005
R3141 DVDD.n457 DVDD.n180 9.3005
R3142 DVDD.n459 DVDD.n458 9.3005
R3143 DVDD.n462 DVDD.n461 9.3005
R3144 DVDD.n463 DVDD.n176 9.3005
R3145 DVDD.n467 DVDD.n466 9.3005
R3146 DVDD.n465 DVDD.n173 9.3005
R3147 DVDD.n472 DVDD.n172 9.3005
R3148 DVDD.n474 DVDD.n473 9.3005
R3149 DVDD.n349 DVDD.n263 9.3005
R3150 DVDD.n353 DVDD.n352 9.3005
R3151 DVDD.n351 DVDD.n260 9.3005
R3152 DVDD.n236 DVDD.n196 9.3005
R3153 DVDD.n190 DVDD.n189 9.3005
R3154 DVDD.n245 DVDD.n244 9.3005
R3155 DVDD.n243 DVDD.n242 9.3005
R3156 DVDD.n366 DVDD.n365 9.3005
R3157 DVDD.n229 DVDD.n228 9.3005
R3158 DVDD.n211 DVDD.n186 9.3005
R3159 DVDD.n208 DVDD.n206 9.3005
R3160 DVDD.n220 DVDD.n219 9.3005
R3161 DVDD.n218 DVDD.n217 9.3005
R3162 DVDD.n213 DVDD.n212 9.3005
R3163 DVDD.n404 DVDD.n403 9.3005
R3164 DVDD.n413 DVDD.n412 9.3005
R3165 DVDD.n410 DVDD.n409 9.3005
R3166 DVDD.n398 DVDD.n397 9.3005
R3167 DVDD.n472 DVDD.n471 9.3005
R3168 DVDD.n468 DVDD.n467 9.3005
R3169 DVDD.n469 DVDD.n173 9.3005
R3170 DVDD.n431 DVDD.n430 9.3005
R3171 DVDD.n433 DVDD.n432 9.3005
R3172 DVDD.n385 DVDD.n382 9.3005
R3173 DVDD.n439 DVDD.n438 9.3005
R3174 DVDD.n441 DVDD.n440 9.3005
R3175 DVDD.n423 DVDD.n422 9.3005
R3176 DVDD.n454 DVDD.n453 9.3005
R3177 DVDD.n341 DVDD.n340 9.3005
R3178 DVDD.n339 DVDD.n265 9.3005
R3179 DVDD.n287 DVDD.n285 9.3005
R3180 DVDD.n289 DVDD.n288 9.3005
R3181 DVDD.n294 DVDD.n293 9.3005
R3182 DVDD.n295 DVDD.n280 9.3005
R3183 DVDD.n297 DVDD.n296 9.3005
R3184 DVDD.n298 DVDD.n279 9.3005
R3185 DVDD.n300 DVDD.n299 9.3005
R3186 DVDD.n301 DVDD.n277 9.3005
R3187 DVDD.n306 DVDD.n275 9.3005
R3188 DVDD.n308 DVDD.n307 9.3005
R3189 DVDD.n309 DVDD.n274 9.3005
R3190 DVDD.n311 DVDD.n310 9.3005
R3191 DVDD.n312 DVDD.n273 9.3005
R3192 DVDD.n314 DVDD.n313 9.3005
R3193 DVDD.n319 DVDD.n269 9.3005
R3194 DVDD.n321 DVDD.n320 9.3005
R3195 DVDD.n329 DVDD.n328 9.3005
R3196 DVDD.n327 DVDD.n325 9.3005
R3197 DVDD.n832 DVDD.n34 9.3005
R3198 DVDD.n834 DVDD.n833 9.3005
R3199 DVDD.n835 DVDD.n33 9.3005
R3200 DVDD.n837 DVDD.n836 9.3005
R3201 DVDD.n839 DVDD.n31 9.3005
R3202 DVDD.n841 DVDD.n840 9.3005
R3203 DVDD.n843 DVDD.n842 9.3005
R3204 DVDD.n844 DVDD.n28 9.3005
R3205 DVDD.n846 DVDD.n845 9.3005
R3206 DVDD.n847 DVDD.n27 9.3005
R3207 DVDD.n849 DVDD.n848 9.3005
R3208 DVDD.n850 DVDD.n26 9.3005
R3209 DVDD.n855 DVDD.n25 9.3005
R3210 DVDD.n857 DVDD.n856 9.3005
R3211 DVDD.n858 DVDD.n24 9.3005
R3212 DVDD.n860 DVDD.n859 9.3005
R3213 DVDD.n862 DVDD.n22 9.3005
R3214 DVDD.n864 DVDD.n863 9.3005
R3215 DVDD.n866 DVDD.n865 9.3005
R3216 DVDD.n867 DVDD.n19 9.3005
R3217 DVDD.n869 DVDD.n868 9.3005
R3218 DVDD.n870 DVDD.n18 9.3005
R3219 DVDD.n872 DVDD.n871 9.3005
R3220 DVDD.n873 DVDD.n17 9.3005
R3221 DVDD.n880 DVDD.n16 9.3005
R3222 DVDD.n882 DVDD.n881 9.3005
R3223 DVDD.n883 DVDD.n15 9.3005
R3224 DVDD.n885 DVDD.n884 9.3005
R3225 DVDD.n886 DVDD.n13 9.3005
R3226 DVDD.n888 DVDD.n887 9.3005
R3227 DVDD.n890 DVDD.n889 9.3005
R3228 DVDD.n891 DVDD.n10 9.3005
R3229 DVDD.n894 DVDD.n893 9.3005
R3230 DVDD.n895 DVDD.n9 9.3005
R3231 DVDD.n897 DVDD.n896 9.3005
R3232 DVDD.n898 DVDD.n8 9.3005
R3233 DVDD.n903 DVDD.n7 9.3005
R3234 DVDD.n905 DVDD.n904 9.3005
R3235 DVDD.n906 DVDD.n6 9.3005
R3236 DVDD.n908 DVDD.n907 9.3005
R3237 DVDD.n909 DVDD.n5 9.3005
R3238 DVDD.n911 DVDD.n910 9.3005
R3239 DVDD.n913 DVDD.n3 9.3005
R3240 DVDD.n917 DVDD.n916 9.3005
R3241 DVDD.n918 DVDD.n2 9.3005
R3242 DVDD.n920 DVDD.n919 9.3005
R3243 DVDD.n921 DVDD.n0 9.3005
R3244 DVDD.n924 DVDD.n923 9.3005
R3245 DVDD.n730 DVDD.n729 9.03579
R3246 DVDD.n763 DVDD.n149 9.03579
R3247 DVDD.n83 DVDD.n73 9.03579
R3248 DVDD.n38 DVDD.n36 9.03579
R3249 DVDD.n724 DVDD.n723 9.03579
R3250 DVDD.n653 DVDD.n646 9.03579
R3251 DVDD.n564 DVDD.n563 9.03579
R3252 DVDD.n582 DVDD.n581 9.03579
R3253 DVDD.n475 DVDD.n474 9.03579
R3254 DVDD.n406 DVDD.n399 9.03579
R3255 DVDD.n248 DVDD.n247 9.03579
R3256 DVDD.n346 DVDD.n345 9.03579
R3257 DVDD.n923 DVDD.n922 9.03579
R3258 DVDD.n899 DVDD.n898 9.03579
R3259 DVDD.n855 DVDD.n854 9.03579
R3260 DVDD.n832 DVDD.n831 9.03579
R3261 DVDD.t176 DVDD.t225 8.879
R3262 DVDD.t254 DVDD.t417 8.879
R3263 DVDD.t165 DVDD.t424 8.879
R3264 DVDD.t247 DVDD.t83 8.879
R3265 DVDD.t126 DVDD.t153 8.879
R3266 DVDD.t474 DVDD.t501 8.879
R3267 DVDD.t113 DVDD.t476 8.879
R3268 DVDD.t131 DVDD.t85 8.879
R3269 DVDD.t19 DVDD.t104 8.879
R3270 DVDD.t340 DVDD.t290 8.879
R3271 DVDD.t226 DVDD.t261 8.879
R3272 DVDD.t237 DVDD.t56 8.879
R3273 DVDD.t440 DVDD.t289 8.879
R3274 DVDD.t23 DVDD.t371 8.879
R3275 DVDD.t401 DVDD.t31 8.879
R3276 DVDD.t172 DVDD.t452 8.879
R3277 DVDD.t342 DVDD.t487 8.879
R3278 DVDD.t514 DVDD.t283 8.879
R3279 DVDD.n477 DVDD.n170 8.86358
R3280 DVDD.n343 DVDD.n342 8.86358
R3281 DVDD.n830 DVDD.n829 8.70378
R3282 DVDD.n727 DVDD.n1 8.70378
R3283 DVDD.n728 DVDD.n727 7.9105
R3284 DVDD.n726 DVDD.n725 7.9105
R3285 DVDD.n477 DVDD.n476 7.9105
R3286 DVDD.n344 DVDD.n343 7.9105
R3287 DVDD.n580 DVDD.n35 7.9105
R3288 DVDD.n829 DVDD.n828 7.9105
R3289 DVDD.n739 DVDD.n161 7.15344
R3290 DVDD.n775 DVDD.n774 7.15344
R3291 DVDD.n95 DVDD.n94 7.15344
R3292 DVDD.n818 DVDD.n47 7.15344
R3293 DVDD.n713 DVDD.n712 7.15344
R3294 DVDD.n665 DVDD.n664 7.15344
R3295 DVDD.n550 DVDD.n513 7.15344
R3296 DVDD.n593 DVDD.n592 7.15344
R3297 DVDD.n464 DVDD.n463 7.15344
R3298 DVDD.n418 DVDD.n417 7.15344
R3299 DVDD.n234 DVDD.n198 7.15344
R3300 DVDD.n357 DVDD.n356 7.15344
R3301 DVDD.n916 DVDD.n915 7.15344
R3302 DVDD.n892 DVDD.n891 7.15344
R3303 DVDD.n862 DVDD.n861 7.15344
R3304 DVDD.n839 DVDD.n838 7.15344
R3305 DVDD.n734 DVDD.n733 6.77697
R3306 DVDD.n760 DVDD.n151 6.77697
R3307 DVDD.n80 DVDD.n79 6.77697
R3308 DVDD.n42 DVDD.n37 6.77697
R3309 DVDD.n720 DVDD.n719 6.77697
R3310 DVDD.n650 DVDD.n648 6.77697
R3311 DVDD.n508 DVDD.n504 6.77697
R3312 DVDD.n586 DVDD.n585 6.77697
R3313 DVDD.n471 DVDD.n470 6.77697
R3314 DVDD.n403 DVDD.n401 6.77697
R3315 DVDD.n193 DVDD.n189 6.77697
R3316 DVDD.n350 DVDD.n349 6.77697
R3317 DVDD.n77 DVDD.n76 6.68889
R3318 DVDD.n758 DVDD.n757 6.68889
R3319 DVDD.n610 DVDD.n609 6.68889
R3320 DVDD.n492 DVDD.n491 6.68889
R3321 DVDD.n374 DVDD.n373 6.68889
R3322 DVDD.n185 DVDD.n184 6.68889
R3323 DVDD.n875 DVDD.n874 6.67829
R3324 DVDD.n852 DVDD.n851 6.67829
R3325 DVDD.n879 DVDD.n878 6.67829
R3326 DVDD.n902 DVDD.n901 6.67829
R3327 DVDD.n742 DVDD.n741 5.64756
R3328 DVDD.n142 DVDD.n137 5.64756
R3329 DVDD.n104 DVDD.n65 5.64756
R3330 DVDD.n816 DVDD.n815 5.64756
R3331 DVDD.n707 DVDD.n485 5.64756
R3332 DVDD.n639 DVDD.n634 5.64756
R3333 DVDD.n548 DVDD.n547 5.64756
R3334 DVDD.n598 DVDD.n572 5.64756
R3335 DVDD.n458 DVDD.n178 5.64756
R3336 DVDD.n392 DVDD.n387 5.64756
R3337 DVDD.n232 DVDD.n231 5.64756
R3338 DVDD.n362 DVDD.n256 5.64756
R3339 DVDD.n912 DVDD.n911 5.64756
R3340 DVDD.n887 DVDD.n12 5.64756
R3341 DVDD.n866 DVDD.n21 5.64756
R3342 DVDD.n843 DVDD.n30 5.64756
R3343 DVDD.n741 DVDD.n740 4.14168
R3344 DVDD.n776 DVDD.n142 4.14168
R3345 DVDD.n96 DVDD.n65 4.14168
R3346 DVDD.n817 DVDD.n816 4.14168
R3347 DVDD.n711 DVDD.n485 4.14168
R3348 DVDD.n666 DVDD.n639 4.14168
R3349 DVDD.n549 DVDD.n548 4.14168
R3350 DVDD.n573 DVDD.n572 4.14168
R3351 DVDD.n462 DVDD.n178 4.14168
R3352 DVDD.n419 DVDD.n392 4.14168
R3353 DVDD.n233 DVDD.n232 4.14168
R3354 DVDD.n257 DVDD.n256 4.14168
R3355 DVDD.n913 DVDD.n912 4.14168
R3356 DVDD.n890 DVDD.n12 4.14168
R3357 DVDD.n863 DVDD.n21 4.14168
R3358 DVDD.n840 DVDD.n30 4.14168
R3359 DVDD.n135 DVDD.n131 3.76521
R3360 DVDD.n111 DVDD.n58 3.76521
R3361 DVDD.n385 DVDD.n381 3.76521
R3362 DVDD.n218 DVDD.n210 3.76521
R3363 DVDD.n163 DVDD.n161 2.63579
R3364 DVDD.n774 DVDD.n772 2.63579
R3365 DVDD.n94 DVDD.n93 2.63579
R3366 DVDD.n47 DVDD.n46 2.63579
R3367 DVDD.n715 DVDD.n713 2.63579
R3368 DVDD.n664 DVDD.n662 2.63579
R3369 DVDD.n555 DVDD.n513 2.63579
R3370 DVDD.n592 DVDD.n591 2.63579
R3371 DVDD.n466 DVDD.n464 2.63579
R3372 DVDD.n417 DVDD.n415 2.63579
R3373 DVDD.n239 DVDD.n198 2.63579
R3374 DVDD.n356 DVDD.n355 2.63579
R3375 DVDD.n915 DVDD.n2 2.63579
R3376 DVDD.n893 DVDD.n892 2.63579
R3377 DVDD.n861 DVDD.n860 2.63579
R3378 DVDD.n838 DVDD.n837 2.63579
R3379 DVDD.n726 DVDD.n477 0.837608
R3380 DVDD.n343 DVDD.n35 0.837608
R3381 DVDD.n328 DVDD.n324 0.753441
R3382 DVDD.n736 DVDD.n166 0.753441
R3383 DVDD.n768 DVDD.n767 0.753441
R3384 DVDD.n89 DVDD.n88 0.753441
R3385 DVDD.n822 DVDD.n821 0.753441
R3386 DVDD.n717 DVDD.n482 0.753441
R3387 DVDD.n658 DVDD.n657 0.753441
R3388 DVDD.n624 DVDD.n497 0.753441
R3389 DVDD.n620 DVDD.n619 0.753441
R3390 DVDD.n559 DVDD.n510 0.753441
R3391 DVDD.n587 DVDD.n575 0.753441
R3392 DVDD.n468 DVDD.n175 0.753441
R3393 DVDD.n411 DVDD.n410 0.753441
R3394 DVDD.n243 DVDD.n195 0.753441
R3395 DVDD.n351 DVDD.n259 0.753441
R3396 DVDD.n319 DVDD.n318 0.753441
R3397 DVDD.n306 DVDD.n305 0.753441
R3398 DVDD.n302 DVDD.n301 0.753441
R3399 DVDD.n288 DVDD.n284 0.753441
R3400 DVDD.n339 DVDD.n338 0.753441
R3401 DVDD.n727 DVDD.n726 0.738527
R3402 DVDD.n829 DVDD.n35 0.738527
R3403 DVDD.n877 DVDD.n876 0.693939
R3404 DVDD.n335 DVDD.n267 0.494563
R3405 DVDD.n332 DVDD.n322 0.494563
R3406 DVDD.n337 DVDD.n336 0.489557
R3407 DVDD.n291 DVDD.n290 0.489557
R3408 DVDD.n317 DVDD.n316 0.489557
R3409 DVDD.n331 DVDD.n330 0.489557
R3410 DVDD.n442 DVDD.n378 0.388044
R3411 DVDD.n292 DVDD.n291 0.387988
R3412 DVDD.n316 DVDD.n315 0.387988
R3413 DVDD.n876 DVDD.n875 0.36602
R3414 DVDD.n878 DVDD.n877 0.36602
R3415 DVDD.n336 DVDD.n335 0.349107
R3416 DVDD.n332 DVDD.n331 0.349107
R3417 DVDD.n853 DVDD.n852 0.305759
R3418 DVDD.n902 DVDD.n900 0.305759
R3419 DVDD.n125 DVDD.n122 0.266946
R3420 DVDD.n304 DVDD.n303 0.21925
R3421 DVDD.n852 DVDD.n26 0.154145
R3422 DVDD.n875 DVDD.n17 0.154145
R3423 DVDD.n878 DVDD.n16 0.154145
R3424 DVDD.n903 DVDD.n902 0.154145
R3425 DVDD.n342 DVDD.n341 0.146169
R3426 DVDD.n285 DVDD.n267 0.146169
R3427 DVDD.n322 DVDD.n321 0.146169
R3428 DVDD.n325 DVDD.n170 0.146169
R3429 DVDD.n337 DVDD.n265 0.141672
R3430 DVDD.n290 DVDD.n289 0.141672
R3431 DVDD.n293 DVDD.n292 0.141672
R3432 DVDD.n315 DVDD.n314 0.141672
R3433 DVDD.n317 DVDD.n269 0.141672
R3434 DVDD.n330 DVDD.n329 0.141672
R3435 DVDD.n78 DVDD.n77 0.136669
R3436 DVDD.n759 DVDD.n758 0.136669
R3437 DVDD.n610 DVDD.n566 0.136669
R3438 DVDD.n649 DVDD.n492 0.136669
R3439 DVDD.n374 DVDD.n250 0.136669
R3440 DVDD.n402 DVDD.n185 0.136669
R3441 DVDD.n122 DVDD.n121 0.136132
R3442 DVDD.n378 DVDD.n186 0.136132
R3443 DVDD.n442 DVDD.n441 0.136132
R3444 DVDD.n622 DVDD.n621 0.122593
R3445 DVDD.n341 DVDD.n265 0.120292
R3446 DVDD.n289 DVDD.n285 0.120292
R3447 DVDD.n293 DVDD.n280 0.120292
R3448 DVDD.n297 DVDD.n280 0.120292
R3449 DVDD.n298 DVDD.n297 0.120292
R3450 DVDD.n299 DVDD.n298 0.120292
R3451 DVDD.n299 DVDD.n277 0.120292
R3452 DVDD.n303 DVDD.n277 0.120292
R3453 DVDD.n304 DVDD.n275 0.120292
R3454 DVDD.n308 DVDD.n275 0.120292
R3455 DVDD.n309 DVDD.n308 0.120292
R3456 DVDD.n310 DVDD.n309 0.120292
R3457 DVDD.n310 DVDD.n273 0.120292
R3458 DVDD.n314 DVDD.n273 0.120292
R3459 DVDD.n321 DVDD.n269 0.120292
R3460 DVDD.n329 DVDD.n325 0.120292
R3461 DVDD.n830 DVDD.n34 0.120292
R3462 DVDD.n834 DVDD.n34 0.120292
R3463 DVDD.n835 DVDD.n834 0.120292
R3464 DVDD.n836 DVDD.n835 0.120292
R3465 DVDD.n836 DVDD.n31 0.120292
R3466 DVDD.n841 DVDD.n31 0.120292
R3467 DVDD.n842 DVDD.n841 0.120292
R3468 DVDD.n842 DVDD.n28 0.120292
R3469 DVDD.n846 DVDD.n28 0.120292
R3470 DVDD.n847 DVDD.n846 0.120292
R3471 DVDD.n848 DVDD.n847 0.120292
R3472 DVDD.n848 DVDD.n26 0.120292
R3473 DVDD.n853 DVDD.n25 0.120292
R3474 DVDD.n857 DVDD.n25 0.120292
R3475 DVDD.n858 DVDD.n857 0.120292
R3476 DVDD.n859 DVDD.n858 0.120292
R3477 DVDD.n859 DVDD.n22 0.120292
R3478 DVDD.n864 DVDD.n22 0.120292
R3479 DVDD.n865 DVDD.n864 0.120292
R3480 DVDD.n865 DVDD.n19 0.120292
R3481 DVDD.n869 DVDD.n19 0.120292
R3482 DVDD.n870 DVDD.n869 0.120292
R3483 DVDD.n871 DVDD.n870 0.120292
R3484 DVDD.n871 DVDD.n17 0.120292
R3485 DVDD.n882 DVDD.n16 0.120292
R3486 DVDD.n883 DVDD.n882 0.120292
R3487 DVDD.n884 DVDD.n883 0.120292
R3488 DVDD.n884 DVDD.n13 0.120292
R3489 DVDD.n888 DVDD.n13 0.120292
R3490 DVDD.n889 DVDD.n888 0.120292
R3491 DVDD.n889 DVDD.n10 0.120292
R3492 DVDD.n894 DVDD.n10 0.120292
R3493 DVDD.n895 DVDD.n894 0.120292
R3494 DVDD.n896 DVDD.n895 0.120292
R3495 DVDD.n896 DVDD.n8 0.120292
R3496 DVDD.n900 DVDD.n8 0.120292
R3497 DVDD.n904 DVDD.n903 0.120292
R3498 DVDD.n904 DVDD.n6 0.120292
R3499 DVDD.n908 DVDD.n6 0.120292
R3500 DVDD.n909 DVDD.n908 0.120292
R3501 DVDD.n910 DVDD.n909 0.120292
R3502 DVDD.n910 DVDD.n3 0.120292
R3503 DVDD.n917 DVDD.n3 0.120292
R3504 DVDD.n918 DVDD.n917 0.120292
R3505 DVDD.n919 DVDD.n918 0.120292
R3506 DVDD.n919 DVDD.n0 0.120292
R3507 DVDD.n924 DVDD.n1 0.120292
R3508 DVDD.n799 DVDD.n798 0.102244
R3509 DVDD DVDD.n0 0.09425
R3510 DVDD.n826 DVDD.n825 0.0673605
R3511 DVDD.n825 DVDD.n824 0.0673605
R3512 DVDD.n824 DVDD.n41 0.0673605
R3513 DVDD.n819 DVDD.n41 0.0673605
R3514 DVDD.n814 DVDD.n44 0.0673605
R3515 DVDD.n807 DVDD.n806 0.0673605
R3516 DVDD.n97 DVDD.n66 0.0673605
R3517 DVDD.n108 DVDD.n62 0.0673605
R3518 DVDD.n126 DVDD.n125 0.0673605
R3519 DVDD.n786 DVDD.n136 0.0673605
R3520 DVDD.n777 DVDD.n141 0.0673605
R3521 DVDD.n751 DVDD.n750 0.0673605
R3522 DVDD.n743 DVDD.n159 0.0673605
R3523 DVDD.n738 DVDD.n737 0.0673605
R3524 DVDD.n737 DVDD.n164 0.0673605
R3525 DVDD.n732 DVDD.n164 0.0673605
R3526 DVDD.n732 DVDD.n731 0.0673605
R3527 DVDD.n583 DVDD.n579 0.0673605
R3528 DVDD.n589 DVDD.n579 0.0673605
R3529 DVDD.n589 DVDD.n576 0.0673605
R3530 DVDD.n594 DVDD.n576 0.0673605
R3531 DVDD.n597 DVDD.n596 0.0673605
R3532 DVDD.n606 DVDD.n605 0.0673605
R3533 DVDD.n551 DVDD.n514 0.0673605
R3534 DVDD.n541 DVDD.n519 0.0673605
R3535 DVDD.n528 DVDD.n526 0.0673605
R3536 DVDD.n621 DVDD.n498 0.0673605
R3537 DVDD.n623 DVDD.n622 0.0673605
R3538 DVDD.n688 DVDD.n495 0.0673605
R3539 DVDD.n676 DVDD.n633 0.0673605
R3540 DVDD.n667 DVDD.n638 0.0673605
R3541 DVDD.n699 DVDD.n698 0.0673605
R3542 DVDD.n710 DVDD.n708 0.0673605
R3543 DVDD.n716 DVDD.n483 0.0673605
R3544 DVDD.n716 DVDD.n480 0.0673605
R3545 DVDD.n721 DVDD.n480 0.0673605
R3546 DVDD.n722 DVDD.n721 0.0673605
R3547 DVDD.n347 DVDD.n263 0.0673605
R3548 DVDD.n353 DVDD.n263 0.0673605
R3549 DVDD.n353 DVDD.n260 0.0673605
R3550 DVDD.n358 DVDD.n260 0.0673605
R3551 DVDD.n361 DVDD.n360 0.0673605
R3552 DVDD.n370 DVDD.n369 0.0673605
R3553 DVDD.n235 DVDD.n199 0.0673605
R3554 DVDD.n225 DVDD.n204 0.0673605
R3555 DVDD.n429 DVDD.n386 0.0673605
R3556 DVDD.n420 DVDD.n391 0.0673605
R3557 DVDD.n450 DVDD.n449 0.0673605
R3558 DVDD.n461 DVDD.n459 0.0673605
R3559 DVDD.n467 DVDD.n176 0.0673605
R3560 DVDD.n467 DVDD.n173 0.0673605
R3561 DVDD.n472 DVDD.n173 0.0673605
R3562 DVDD.n473 DVDD.n472 0.0673605
R3563 DVDD.n162 DVDD.n159 0.056111
R3564 DVDD.n728 DVDD.n167 0.056111
R3565 DVDD.n828 DVDD.n827 0.056111
R3566 DVDD.n820 DVDD.n44 0.056111
R3567 DVDD.n710 DVDD.n709 0.056111
R3568 DVDD.n725 DVDD.n478 0.056111
R3569 DVDD.n584 DVDD.n580 0.056111
R3570 DVDD.n596 DVDD.n595 0.056111
R3571 DVDD.n461 DVDD.n460 0.056111
R3572 DVDD.n476 DVDD.n171 0.056111
R3573 DVDD.n348 DVDD.n344 0.056111
R3574 DVDD.n360 DVDD.n359 0.056111
R3575 DVDD.n814 DVDD.n813 0.0557326
R3576 DVDD.n811 DVDD.n50 0.0557326
R3577 DVDD.n810 DVDD.n52 0.0557326
R3578 DVDD.n747 DVDD.n154 0.0557326
R3579 DVDD.n746 DVDD.n157 0.0557326
R3580 DVDD.n744 DVDD.n743 0.0557326
R3581 DVDD.n597 DVDD.n569 0.0557326
R3582 DVDD.n601 DVDD.n600 0.0557326
R3583 DVDD.n604 DVDD.n568 0.0557326
R3584 DVDD.n704 DVDD.n700 0.0557326
R3585 DVDD.n703 DVDD.n487 0.0557326
R3586 DVDD.n708 DVDD.n486 0.0557326
R3587 DVDD.n361 DVDD.n253 0.0557326
R3588 DVDD.n365 DVDD.n364 0.0557326
R3589 DVDD.n368 DVDD.n252 0.0557326
R3590 DVDD.n455 DVDD.n451 0.0557326
R3591 DVDD.n454 DVDD.n180 0.0557326
R3592 DVDD.n459 DVDD.n179 0.0557326
R3593 DVDD.n109 DVDD.n61 0.0470116
R3594 DVDD.n114 DVDD.n113 0.0470116
R3595 DVDD.n117 DVDD.n59 0.0470116
R3596 DVDD.n118 DVDD.n56 0.0470116
R3597 DVDD.n128 DVDD.n123 0.0470116
R3598 DVDD.n795 DVDD.n129 0.0470116
R3599 DVDD.n794 DVDD.n132 0.0470116
R3600 DVDD.n791 DVDD.n790 0.0470116
R3601 DVDD.n787 DVDD.n134 0.0470116
R3602 DVDD.n537 DVDD.n521 0.0470116
R3603 DVDD.n536 DVDD.n522 0.0470116
R3604 DVDD.n532 DVDD.n531 0.0470116
R3605 DVDD.n529 DVDD.n525 0.0470116
R3606 DVDD.n684 DVDD.n627 0.0470116
R3607 DVDD.n683 DVDD.n628 0.0470116
R3608 DVDD.n680 DVDD.n679 0.0470116
R3609 DVDD.n677 DVDD.n630 0.0470116
R3610 DVDD.n221 DVDD.n206 0.0470116
R3611 DVDD.n220 DVDD.n207 0.0470116
R3612 DVDD.n217 DVDD.n216 0.0470116
R3613 DVDD.n214 DVDD.n213 0.0470116
R3614 DVDD.n438 DVDD.n379 0.0470116
R3615 DVDD.n437 DVDD.n382 0.0470116
R3616 DVDD.n434 DVDD.n433 0.0470116
R3617 DVDD.n430 DVDD.n384 0.0470116
R3618 DVDD.n806 DVDD.n805 0.0441047
R3619 DVDD.n55 DVDD.n54 0.0441047
R3620 DVDD.n81 DVDD.n74 0.0441047
R3621 DVDD.n82 DVDD.n72 0.0441047
R3622 DVDD.n87 DVDD.n85 0.0441047
R3623 DVDD.n86 DVDD.n69 0.0441047
R3624 DVDD.n92 DVDD.n91 0.0441047
R3625 DVDD.n771 DVDD.n144 0.0441047
R3626 DVDD.n770 DVDD.n145 0.0441047
R3627 DVDD.n766 DVDD.n765 0.0441047
R3628 DVDD.n762 DVDD.n148 0.0441047
R3629 DVDD.n761 DVDD.n150 0.0441047
R3630 DVDD.n755 DVDD.n152 0.0441047
R3631 DVDD.n754 DVDD.n751 0.0441047
R3632 DVDD.n606 DVDD.n502 0.0441047
R3633 DVDD.n611 DVDD.n503 0.0441047
R3634 DVDD.n565 DVDD.n505 0.0441047
R3635 DVDD.n562 DVDD.n561 0.0441047
R3636 DVDD.n558 DVDD.n507 0.0441047
R3637 DVDD.n557 DVDD.n511 0.0441047
R3638 DVDD.n554 DVDD.n553 0.0441047
R3639 DVDD.n661 DVDD.n641 0.0441047
R3640 DVDD.n660 DVDD.n642 0.0441047
R3641 DVDD.n656 DVDD.n655 0.0441047
R3642 DVDD.n652 DVDD.n645 0.0441047
R3643 DVDD.n651 DVDD.n647 0.0441047
R3644 DVDD.n695 DVDD.n694 0.0441047
R3645 DVDD.n698 DVDD.n490 0.0441047
R3646 DVDD.n370 DVDD.n187 0.0441047
R3647 DVDD.n375 DVDD.n188 0.0441047
R3648 DVDD.n249 DVDD.n190 0.0441047
R3649 DVDD.n246 DVDD.n245 0.0441047
R3650 DVDD.n242 DVDD.n192 0.0441047
R3651 DVDD.n241 DVDD.n196 0.0441047
R3652 DVDD.n238 DVDD.n237 0.0441047
R3653 DVDD.n414 DVDD.n394 0.0441047
R3654 DVDD.n413 DVDD.n395 0.0441047
R3655 DVDD.n409 DVDD.n408 0.0441047
R3656 DVDD.n405 DVDD.n398 0.0441047
R3657 DVDD.n404 DVDD.n400 0.0441047
R3658 DVDD.n446 DVDD.n445 0.0441047
R3659 DVDD.n449 DVDD.n183 0.0441047
R3660 DVDD.n77 DVDD.n55 0.042901
R3661 DVDD.n758 DVDD.n152 0.042901
R3662 DVDD.n611 DVDD.n610 0.042901
R3663 DVDD.n694 DVDD.n492 0.042901
R3664 DVDD.n375 DVDD.n374 0.042901
R3665 DVDD.n445 DVDD.n185 0.042901
R3666 DVDD.n78 DVDD.n74 0.0359214
R3667 DVDD.n759 DVDD.n150 0.0359214
R3668 DVDD.n566 DVDD.n565 0.0359214
R3669 DVDD.n649 DVDD.n647 0.0359214
R3670 DVDD.n250 DVDD.n249 0.0359214
R3671 DVDD.n402 DVDD.n400 0.0359214
R3672 DVDD.n103 DVDD.n98 0.0353837
R3673 DVDD.n102 DVDD.n63 0.0353837
R3674 DVDD.n99 DVDD.n62 0.0353837
R3675 DVDD.n138 DVDD.n136 0.0353837
R3676 DVDD.n781 DVDD.n780 0.0353837
R3677 DVDD.n778 DVDD.n139 0.0353837
R3678 DVDD.n546 DVDD.n517 0.0353837
R3679 DVDD.n545 DVDD.n518 0.0353837
R3680 DVDD.n542 DVDD.n541 0.0353837
R3681 DVDD.n526 DVDD.n501 0.0353837
R3682 DVDD.n617 DVDD.n616 0.0353837
R3683 DVDD.n494 DVDD.n493 0.0353837
R3684 DVDD.n689 DVDD.n688 0.0353837
R3685 DVDD.n635 DVDD.n633 0.0353837
R3686 DVDD.n671 DVDD.n670 0.0353837
R3687 DVDD.n668 DVDD.n636 0.0353837
R3688 DVDD.n230 DVDD.n202 0.0353837
R3689 DVDD.n229 DVDD.n203 0.0353837
R3690 DVDD.n226 DVDD.n225 0.0353837
R3691 DVDD.n388 DVDD.n386 0.0353837
R3692 DVDD.n424 DVDD.n423 0.0353837
R3693 DVDD.n421 DVDD.n389 0.0353837
R3694 DVDD.n98 DVDD.n97 0.0324767
R3695 DVDD.n103 DVDD.n102 0.0324767
R3696 DVDD.n99 DVDD.n63 0.0324767
R3697 DVDD.n781 DVDD.n138 0.0324767
R3698 DVDD.n780 DVDD.n139 0.0324767
R3699 DVDD.n778 DVDD.n777 0.0324767
R3700 DVDD.n517 DVDD.n514 0.0324767
R3701 DVDD.n546 DVDD.n545 0.0324767
R3702 DVDD.n542 DVDD.n518 0.0324767
R3703 DVDD.n617 DVDD.n501 0.0324767
R3704 DVDD.n616 DVDD.n498 0.0324767
R3705 DVDD.n623 DVDD.n493 0.0324767
R3706 DVDD.n689 DVDD.n494 0.0324767
R3707 DVDD.n671 DVDD.n635 0.0324767
R3708 DVDD.n670 DVDD.n636 0.0324767
R3709 DVDD.n668 DVDD.n667 0.0324767
R3710 DVDD.n202 DVDD.n199 0.0324767
R3711 DVDD.n230 DVDD.n229 0.0324767
R3712 DVDD.n226 DVDD.n203 0.0324767
R3713 DVDD.n424 DVDD.n388 0.0324767
R3714 DVDD.n423 DVDD.n389 0.0324767
R3715 DVDD.n421 DVDD.n420 0.0324767
R3716 DVDD DVDD.n924 0.0265417
R3717 DVDD.n805 DVDD.n54 0.0237558
R3718 DVDD.n82 DVDD.n81 0.0237558
R3719 DVDD.n85 DVDD.n72 0.0237558
R3720 DVDD.n87 DVDD.n86 0.0237558
R3721 DVDD.n92 DVDD.n69 0.0237558
R3722 DVDD.n91 DVDD.n66 0.0237558
R3723 DVDD.n144 DVDD.n141 0.0237558
R3724 DVDD.n771 DVDD.n770 0.0237558
R3725 DVDD.n766 DVDD.n145 0.0237558
R3726 DVDD.n765 DVDD.n148 0.0237558
R3727 DVDD.n762 DVDD.n761 0.0237558
R3728 DVDD.n755 DVDD.n754 0.0237558
R3729 DVDD.n503 DVDD.n502 0.0237558
R3730 DVDD.n562 DVDD.n505 0.0237558
R3731 DVDD.n561 DVDD.n507 0.0237558
R3732 DVDD.n558 DVDD.n557 0.0237558
R3733 DVDD.n554 DVDD.n511 0.0237558
R3734 DVDD.n553 DVDD.n551 0.0237558
R3735 DVDD.n641 DVDD.n638 0.0237558
R3736 DVDD.n661 DVDD.n660 0.0237558
R3737 DVDD.n656 DVDD.n642 0.0237558
R3738 DVDD.n655 DVDD.n645 0.0237558
R3739 DVDD.n652 DVDD.n651 0.0237558
R3740 DVDD.n695 DVDD.n490 0.0237558
R3741 DVDD.n188 DVDD.n187 0.0237558
R3742 DVDD.n246 DVDD.n190 0.0237558
R3743 DVDD.n245 DVDD.n192 0.0237558
R3744 DVDD.n242 DVDD.n241 0.0237558
R3745 DVDD.n238 DVDD.n196 0.0237558
R3746 DVDD.n237 DVDD.n235 0.0237558
R3747 DVDD.n394 DVDD.n391 0.0237558
R3748 DVDD.n414 DVDD.n413 0.0237558
R3749 DVDD.n409 DVDD.n395 0.0237558
R3750 DVDD.n408 DVDD.n398 0.0237558
R3751 DVDD.n405 DVDD.n404 0.0237558
R3752 DVDD.n446 DVDD.n183 0.0237558
R3753 DVDD.n109 DVDD.n108 0.0208488
R3754 DVDD.n113 DVDD.n61 0.0208488
R3755 DVDD.n114 DVDD.n59 0.0208488
R3756 DVDD.n118 DVDD.n117 0.0208488
R3757 DVDD.n121 DVDD.n56 0.0208488
R3758 DVDD.n126 DVDD.n123 0.0208488
R3759 DVDD.n799 DVDD.n128 0.0208488
R3760 DVDD.n798 DVDD.n129 0.0208488
R3761 DVDD.n795 DVDD.n794 0.0208488
R3762 DVDD.n791 DVDD.n132 0.0208488
R3763 DVDD.n790 DVDD.n134 0.0208488
R3764 DVDD.n787 DVDD.n786 0.0208488
R3765 DVDD.n521 DVDD.n519 0.0208488
R3766 DVDD.n537 DVDD.n536 0.0208488
R3767 DVDD.n532 DVDD.n522 0.0208488
R3768 DVDD.n531 DVDD.n525 0.0208488
R3769 DVDD.n529 DVDD.n528 0.0208488
R3770 DVDD.n627 DVDD.n495 0.0208488
R3771 DVDD.n684 DVDD.n683 0.0208488
R3772 DVDD.n680 DVDD.n628 0.0208488
R3773 DVDD.n679 DVDD.n630 0.0208488
R3774 DVDD.n677 DVDD.n676 0.0208488
R3775 DVDD.n206 DVDD.n204 0.0208488
R3776 DVDD.n221 DVDD.n220 0.0208488
R3777 DVDD.n217 DVDD.n207 0.0208488
R3778 DVDD.n216 DVDD.n213 0.0208488
R3779 DVDD.n214 DVDD.n186 0.0208488
R3780 DVDD.n441 DVDD.n379 0.0208488
R3781 DVDD.n438 DVDD.n437 0.0208488
R3782 DVDD.n434 DVDD.n382 0.0208488
R3783 DVDD.n433 DVDD.n384 0.0208488
R3784 DVDD.n430 DVDD.n429 0.0208488
R3785 DVDD.n827 DVDD.n826 0.0126656
R3786 DVDD.n820 DVDD.n819 0.0126656
R3787 DVDD.n738 DVDD.n162 0.0126656
R3788 DVDD.n731 DVDD.n167 0.0126656
R3789 DVDD.n584 DVDD.n583 0.0126656
R3790 DVDD.n595 DVDD.n594 0.0126656
R3791 DVDD.n709 DVDD.n483 0.0126656
R3792 DVDD.n722 DVDD.n478 0.0126656
R3793 DVDD.n348 DVDD.n347 0.0126656
R3794 DVDD.n359 DVDD.n358 0.0126656
R3795 DVDD.n460 DVDD.n176 0.0126656
R3796 DVDD.n473 DVDD.n171 0.0126656
R3797 DVDD.n813 DVDD.n50 0.0121279
R3798 DVDD.n811 DVDD.n810 0.0121279
R3799 DVDD.n807 DVDD.n52 0.0121279
R3800 DVDD.n750 DVDD.n154 0.0121279
R3801 DVDD.n747 DVDD.n746 0.0121279
R3802 DVDD.n744 DVDD.n157 0.0121279
R3803 DVDD.n600 DVDD.n569 0.0121279
R3804 DVDD.n601 DVDD.n568 0.0121279
R3805 DVDD.n605 DVDD.n604 0.0121279
R3806 DVDD.n700 DVDD.n699 0.0121279
R3807 DVDD.n704 DVDD.n703 0.0121279
R3808 DVDD.n487 DVDD.n486 0.0121279
R3809 DVDD.n364 DVDD.n253 0.0121279
R3810 DVDD.n365 DVDD.n252 0.0121279
R3811 DVDD.n369 DVDD.n368 0.0121279
R3812 DVDD.n451 DVDD.n450 0.0121279
R3813 DVDD.n455 DVDD.n454 0.0121279
R3814 DVDD.n180 DVDD.n179 0.0121279
R3815 A15.n1 A15.t8 373.283
R3816 A15.n0 A15.t10 347.577
R3817 A15.n9 A15.t4 334.723
R3818 A15.n3 A15.t5 323.476
R3819 A15.n3 A15.t11 217.436
R3820 A15.n5 A15.t1 212.081
R3821 A15.n6 A15.t3 212.081
R3822 A15.n9 A15.t6 206.19
R3823 A15.n0 A15.t9 193.337
R3824 A15.n8 A15.n7 174.552
R3825 A15.n4 A15.n3 169.833
R3826 A15.n1 A15.t7 167.63
R3827 A15.n2 A15.n0 166.843
R3828 A15.n2 A15.n1 166.421
R3829 A15.n10 A15.n9 152
R3830 A15.n5 A15.t0 139.78
R3831 A15.n6 A15.t2 139.78
R3832 A15.n7 A15.n5 37.246
R3833 A15.n7 A15.n6 24.1005
R3834 A15.n10 A15.n8 17.5294
R3835 A15.n4 A15.n2 1.55989
R3836 A15 A15.n10 0.914786
R3837 A15.n8 A15.n4 0.112749
R3838 A2.n1 A2.t0 373.283
R3839 A2.n0 A2.t11 347.577
R3840 A2.n9 A2.t4 334.723
R3841 A2.n3 A2.t3 323.476
R3842 A2.n3 A2.t6 217.436
R3843 A2.n5 A2.t8 212.081
R3844 A2.n6 A2.t1 212.081
R3845 A2.n9 A2.t2 206.19
R3846 A2.n0 A2.t9 193.337
R3847 A2.n8 A2.n7 171.9
R3848 A2.n4 A2.n3 169.833
R3849 A2.n1 A2.t5 167.63
R3850 A2.n2 A2.n0 166.843
R3851 A2.n2 A2.n1 166.421
R3852 A2.n10 A2.n9 152
R3853 A2.n5 A2.t7 139.78
R3854 A2.n6 A2.t10 139.78
R3855 A2.n7 A2.n6 37.246
R3856 A2.n7 A2.n5 24.1005
R3857 A2.n10 A2.n8 17.5294
R3858 A2 A2.n10 2.74336
R3859 A2.n4 A2.n2 1.55989
R3860 A2.n8 A2.n4 0.112749
R3861 B14.n9 B14.t9 384.529
R3862 B14.n3 B14.t3 373.283
R3863 B14.n5 B14.t5 351.861
R3864 B14.n4 B14.t10 297.233
R3865 B14.n2 B14.n1 263.558
R3866 B14.n0 B14.t6 241.536
R3867 B14.n1 B14.t8 241.536
R3868 B14.n6 B14.n5 214.362
R3869 B14.n0 B14.t4 169.237
R3870 B14.n1 B14.t7 169.237
R3871 B14.n7 B14.n3 167.825
R3872 B14.n3 B14.t0 167.63
R3873 B14.n7 B14.n6 163.79
R3874 B14.n9 B14.t1 156.382
R3875 B14.n2 B14.n0 152.298
R3876 B14.n10 B14.n9 152
R3877 B14.n5 B14.t11 109.215
R3878 B14.n4 B14.t2 102.659
R3879 B14.n6 B14.n4 47.4474
R3880 B14.n8 B14.n2 19.8357
R3881 B14.n10 B14.n8 16.0683
R3882 B14.n8 B14.n7 1.54462
R3883 B14 B14.n10 0.589006
R3884 B9.n0 B9.t1 384.529
R3885 B9.n4 B9.t10 373.283
R3886 B9.n6 B9.t0 351.861
R3887 B9.n5 B9.t7 297.233
R3888 B9.n3 B9.n2 257.209
R3889 B9.n1 B9.t6 241.536
R3890 B9.n2 B9.t2 241.536
R3891 B9.n7 B9.n6 214.362
R3892 B9.n1 B9.t3 169.237
R3893 B9.n2 B9.t9 169.237
R3894 B9.n8 B9.n4 167.825
R3895 B9.n4 B9.t4 167.63
R3896 B9.n8 B9.n7 163.79
R3897 B9.n0 B9.t8 156.382
R3898 B9.n3 B9.n1 153.97
R3899 B9 B9.n0 152.883
R3900 B9.n6 B9.t5 109.215
R3901 B9.n5 B9.t11 102.659
R3902 B9.n7 B9.n5 47.4474
R3903 B9.n9 B9.n3 20.0296
R3904 B9 B9.n9 15.1856
R3905 B9.n9 B9.n8 1.54462
R3906 A10.n1 A10.t4 373.283
R3907 A10.n0 A10.t5 347.577
R3908 A10.n9 A10.t3 334.723
R3909 A10.n3 A10.t11 323.476
R3910 A10.n3 A10.t7 217.436
R3911 A10.n5 A10.t8 212.081
R3912 A10.n6 A10.t2 212.081
R3913 A10.n9 A10.t10 206.19
R3914 A10.n0 A10.t1 193.337
R3915 A10.n8 A10.n7 171.9
R3916 A10.n4 A10.n3 169.833
R3917 A10.n1 A10.t0 167.63
R3918 A10.n2 A10.n0 166.843
R3919 A10.n2 A10.n1 166.421
R3920 A10.n10 A10.n9 152
R3921 A10.n5 A10.t6 139.78
R3922 A10.n6 A10.t9 139.78
R3923 A10.n7 A10.n5 37.246
R3924 A10.n7 A10.n6 24.1005
R3925 A10.n10 A10.n8 17.5294
R3926 A10 A10.n10 2.74336
R3927 A10.n4 A10.n2 1.55989
R3928 A10.n8 A10.n4 0.112749
R3929 A14.n1 A14.t3 373.283
R3930 A14.n0 A14.t7 347.577
R3931 A14.n9 A14.t5 334.723
R3932 A14.n3 A14.t2 323.476
R3933 A14.n3 A14.t8 217.436
R3934 A14.n5 A14.t6 212.081
R3935 A14.n6 A14.t10 212.081
R3936 A14.n9 A14.t11 206.19
R3937 A14.n0 A14.t1 193.337
R3938 A14.n8 A14.n7 171.9
R3939 A14.n4 A14.n3 169.833
R3940 A14.n1 A14.t0 167.63
R3941 A14.n2 A14.n0 166.843
R3942 A14.n2 A14.n1 166.421
R3943 A14.n10 A14.n9 152
R3944 A14.n5 A14.t4 139.78
R3945 A14.n6 A14.t9 139.78
R3946 A14.n7 A14.n5 37.246
R3947 A14.n7 A14.n6 24.1005
R3948 A14.n10 A14.n8 17.5294
R3949 A14 A14.n10 2.74336
R3950 A14.n4 A14.n2 1.55989
R3951 A14.n8 A14.n4 0.112749
R3952 A1.n1 A1.t3 373.283
R3953 A1.n0 A1.t10 347.577
R3954 A1.n9 A1.t1 334.723
R3955 A1.n3 A1.t9 323.476
R3956 A1.n3 A1.t8 217.436
R3957 A1.n5 A1.t11 212.081
R3958 A1.n6 A1.t4 212.081
R3959 A1.n9 A1.t0 206.19
R3960 A1.n0 A1.t6 193.337
R3961 A1.n8 A1.n7 174.552
R3962 A1.n4 A1.n3 169.833
R3963 A1.n1 A1.t5 167.63
R3964 A1.n2 A1.n0 166.843
R3965 A1.n2 A1.n1 166.421
R3966 A1.n10 A1.n9 152
R3967 A1.n5 A1.t7 139.78
R3968 A1.n6 A1.t2 139.78
R3969 A1.n7 A1.n6 37.246
R3970 A1.n7 A1.n5 24.1005
R3971 A1.n10 A1.n8 17.5294
R3972 A1 A1.n10 3.2005
R3973 A1.n4 A1.n2 1.55989
R3974 A1.n8 A1.n4 0.112749
R3975 A6.n1 A6.t7 373.283
R3976 A6.n0 A6.t3 347.577
R3977 A6.n9 A6.t4 334.723
R3978 A6.n3 A6.t0 323.476
R3979 A6.n3 A6.t8 217.436
R3980 A6.n5 A6.t2 212.081
R3981 A6.n6 A6.t5 212.081
R3982 A6.n9 A6.t1 206.19
R3983 A6.n0 A6.t10 193.337
R3984 A6.n8 A6.n7 171.9
R3985 A6.n4 A6.n3 169.833
R3986 A6.n1 A6.t6 167.63
R3987 A6.n2 A6.n0 166.843
R3988 A6.n2 A6.n1 166.421
R3989 A6.n10 A6.n9 152
R3990 A6.n5 A6.t9 139.78
R3991 A6.n6 A6.t11 139.78
R3992 A6.n7 A6.n6 37.246
R3993 A6.n7 A6.n5 24.1005
R3994 A6.n10 A6.n8 17.5294
R3995 A6 A6.n10 2.74336
R3996 A6.n4 A6.n2 1.55989
R3997 A6.n8 A6.n4 0.112749
R3998 A8.n1 A8.t3 373.283
R3999 A8.n0 A8.t4 347.577
R4000 A8.n9 A8.t1 334.723
R4001 A8.n3 A8.t0 323.476
R4002 A8.n3 A8.t5 217.436
R4003 A8.n5 A8.t6 212.081
R4004 A8.n6 A8.t11 212.081
R4005 A8.n9 A8.t8 206.19
R4006 A8.n0 A8.t10 193.337
R4007 A8.n8 A8.n7 171.9
R4008 A8.n4 A8.n3 169.833
R4009 A8.n1 A8.t9 167.63
R4010 A8.n2 A8.n0 166.843
R4011 A8.n2 A8.n1 166.421
R4012 A8.n10 A8.n9 152
R4013 A8.n5 A8.t2 139.78
R4014 A8.n6 A8.t7 139.78
R4015 A8.n7 A8.n5 37.246
R4016 A8.n7 A8.n6 24.1005
R4017 A8.n10 A8.n8 17.5294
R4018 A8 A8.n10 2.05764
R4019 A8.n4 A8.n2 1.55989
R4020 A8.n8 A8.n4 0.112749
R4021 B2.n9 B2.t11 384.529
R4022 B2.n0 B2.t2 373.283
R4023 B2.n2 B2.t9 351.861
R4024 B2.n1 B2.t10 297.233
R4025 B2.n7 B2.n5 263.558
R4026 B2.n6 B2.t3 241.536
R4027 B2.n5 B2.t4 241.536
R4028 B2.n3 B2.n2 214.362
R4029 B2.n6 B2.t0 169.237
R4030 B2.n5 B2.t1 169.237
R4031 B2.n4 B2.n0 167.825
R4032 B2.n0 B2.t7 167.63
R4033 B2.n4 B2.n3 163.79
R4034 B2.n9 B2.t6 156.382
R4035 B2.n7 B2.n6 152.298
R4036 B2.n10 B2.n9 152
R4037 B2.n2 B2.t8 109.215
R4038 B2.n1 B2.t5 102.659
R4039 B2.n3 B2.n1 47.4474
R4040 B2.n8 B2.n7 19.8357
R4041 B2.n10 B2.n8 16.0683
R4042 B2.n8 B2.n4 1.54462
R4043 B2 B2.n10 0.589006
R4044 B6.n9 B6.t9 384.529
R4045 B6.n0 B6.t2 373.283
R4046 B6.n2 B6.t8 351.861
R4047 B6.n1 B6.t10 297.233
R4048 B6.n7 B6.n5 263.558
R4049 B6.n6 B6.t4 241.536
R4050 B6.n5 B6.t5 241.536
R4051 B6.n3 B6.n2 214.362
R4052 B6.n6 B6.t0 169.237
R4053 B6.n5 B6.t1 169.237
R4054 B6.n4 B6.n0 167.825
R4055 B6.n0 B6.t3 167.63
R4056 B6.n4 B6.n3 163.79
R4057 B6.n9 B6.t11 156.382
R4058 B6.n7 B6.n6 152.298
R4059 B6.n10 B6.n9 152
R4060 B6.n2 B6.t6 109.215
R4061 B6.n1 B6.t7 102.659
R4062 B6.n3 B6.n1 47.4474
R4063 B6.n8 B6.n7 19.8357
R4064 B6.n10 B6.n8 16.0683
R4065 B6.n8 B6.n4 1.54462
R4066 B6 B6.n10 0.589006
R4067 A4.n1 A4.t8 373.283
R4068 A4.n0 A4.t3 347.577
R4069 A4.n9 A4.t5 334.723
R4070 A4.n3 A4.t1 323.476
R4071 A4.n3 A4.t6 217.436
R4072 A4.n5 A4.t0 212.081
R4073 A4.n6 A4.t2 212.081
R4074 A4.n9 A4.t11 206.19
R4075 A4.n0 A4.t9 193.337
R4076 A4.n8 A4.n7 171.9
R4077 A4.n4 A4.n3 169.833
R4078 A4.n1 A4.t4 167.63
R4079 A4.n2 A4.n0 166.843
R4080 A4.n2 A4.n1 166.421
R4081 A4.n10 A4.n9 152
R4082 A4.n5 A4.t7 139.78
R4083 A4.n6 A4.t10 139.78
R4084 A4.n7 A4.n6 37.246
R4085 A4.n7 A4.n5 24.1005
R4086 A4.n10 A4.n8 17.5294
R4087 A4 A4.n10 2.28621
R4088 A4.n4 A4.n2 1.55989
R4089 A4.n8 A4.n4 0.112749
R4090 B13.n0 B13.t2 384.529
R4091 B13.n4 B13.t0 373.283
R4092 B13.n6 B13.t10 351.861
R4093 B13.n5 B13.t7 297.233
R4094 B13.n3 B13.n2 257.209
R4095 B13.n1 B13.t11 241.536
R4096 B13.n2 B13.t9 241.536
R4097 B13.n7 B13.n6 214.362
R4098 B13.n1 B13.t8 169.237
R4099 B13.n2 B13.t6 169.237
R4100 B13.n8 B13.n4 167.825
R4101 B13.n4 B13.t4 167.63
R4102 B13.n8 B13.n7 163.79
R4103 B13.n0 B13.t1 156.382
R4104 B13.n3 B13.n1 153.97
R4105 B13 B13.n0 152.294
R4106 B13.n6 B13.t5 109.215
R4107 B13.n5 B13.t3 102.659
R4108 B13.n7 B13.n5 47.4474
R4109 B13.n9 B13.n3 20.0296
R4110 B13 B13.n9 15.7741
R4111 B13.n9 B13.n8 1.54462
R4112 B10.n9 B10.t6 384.529
R4113 B10.n3 B10.t1 373.283
R4114 B10.n5 B10.t3 351.861
R4115 B10.n4 B10.t7 297.233
R4116 B10.n2 B10.n1 263.558
R4117 B10.n0 B10.t8 241.536
R4118 B10.n1 B10.t10 241.536
R4119 B10.n6 B10.n5 214.362
R4120 B10.n0 B10.t2 169.237
R4121 B10.n1 B10.t4 169.237
R4122 B10.n7 B10.n3 167.825
R4123 B10.n3 B10.t5 167.63
R4124 B10.n7 B10.n6 163.79
R4125 B10.n9 B10.t11 156.382
R4126 B10.n2 B10.n0 152.298
R4127 B10.n10 B10.n9 152
R4128 B10.n5 B10.t9 109.215
R4129 B10.n4 B10.t0 102.659
R4130 B10.n6 B10.n4 47.4474
R4131 B10.n8 B10.n2 19.8357
R4132 B10.n10 B10.n8 16.0683
R4133 B10.n8 B10.n7 1.54462
R4134 B10 B10.n10 0.589006
R4135 A13.n1 A13.t8 373.283
R4136 A13.n0 A13.t6 347.577
R4137 A13.n9 A13.t1 334.723
R4138 A13.n3 A13.t4 323.476
R4139 A13.n3 A13.t2 217.436
R4140 A13.n5 A13.t9 212.081
R4141 A13.n6 A13.t0 212.081
R4142 A13.n9 A13.t10 206.19
R4143 A13.n0 A13.t3 193.337
R4144 A13.n8 A13.n7 174.552
R4145 A13.n4 A13.n3 169.833
R4146 A13.n1 A13.t7 167.63
R4147 A13.n2 A13.n0 166.843
R4148 A13.n2 A13.n1 166.421
R4149 A13.n10 A13.n9 152
R4150 A13.n5 A13.t5 139.78
R4151 A13.n6 A13.t11 139.78
R4152 A13.n7 A13.n5 37.246
R4153 A13.n7 A13.n6 24.1005
R4154 A13.n10 A13.n8 17.5294
R4155 A13 A13.n10 3.2005
R4156 A13.n4 A13.n2 1.55989
R4157 A13.n8 A13.n4 0.112749
R4158 B0.n9 B0.t10 384.529
R4159 B0.n0 B0.t4 373.283
R4160 B0.n2 B0.t9 351.861
R4161 B0.n1 B0.t11 297.233
R4162 B0.n7 B0.n5 263.558
R4163 B0.n6 B0.t6 241.536
R4164 B0.n5 B0.t0 241.536
R4165 B0.n3 B0.n2 214.362
R4166 B0.n6 B0.t3 169.237
R4167 B0.n5 B0.t8 169.237
R4168 B0.n4 B0.n0 167.825
R4169 B0.n0 B0.t5 167.63
R4170 B0.n4 B0.n3 163.79
R4171 B0.n9 B0.t7 156.382
R4172 B0 B0.n9 154.649
R4173 B0.n7 B0.n6 152.298
R4174 B0.n2 B0.t2 109.215
R4175 B0.n1 B0.t1 102.659
R4176 B0.n3 B0.n1 47.4474
R4177 B0.n8 B0.n7 19.8357
R4178 B0 B0.n8 13.42
R4179 B0.n8 B0.n4 1.54462
R4180 A7.n1 A7.t2 373.283
R4181 A7.n0 A7.t10 347.577
R4182 A7.n9 A7.t5 334.723
R4183 A7.n3 A7.t4 323.476
R4184 A7.n3 A7.t0 217.436
R4185 A7.n5 A7.t9 212.081
R4186 A7.n6 A7.t8 212.081
R4187 A7.n9 A7.t1 206.19
R4188 A7.n0 A7.t7 193.337
R4189 A7.n8 A7.n7 174.552
R4190 A7.n4 A7.n3 169.833
R4191 A7.n1 A7.t11 167.63
R4192 A7.n2 A7.n0 166.843
R4193 A7.n2 A7.n1 166.421
R4194 A7.n10 A7.n9 152
R4195 A7.n5 A7.t6 139.78
R4196 A7.n6 A7.t3 139.78
R4197 A7.n7 A7.n6 37.246
R4198 A7.n7 A7.n5 24.1005
R4199 A7.n10 A7.n8 17.5294
R4200 A7.n10 A7 14.0805
R4201 A7 A7.n10 2.51479
R4202 A7.n4 A7.n2 1.55989
R4203 A7.n8 A7.n4 0.112749
R4204 B8.n0 B8.t6 384.529
R4205 B8.n4 B8.t2 373.283
R4206 B8.n6 B8.t4 351.861
R4207 B8.n5 B8.t11 297.233
R4208 B8.n3 B8.n2 263.558
R4209 B8.n1 B8.t7 241.536
R4210 B8.n2 B8.t9 241.536
R4211 B8.n7 B8.n6 214.362
R4212 B8.n1 B8.t3 169.237
R4213 B8.n2 B8.t5 169.237
R4214 B8.n8 B8.n4 167.825
R4215 B8.n4 B8.t10 167.63
R4216 B8.n8 B8.n7 163.79
R4217 B8.n0 B8.t0 156.382
R4218 B8 B8.n0 152.441
R4219 B8.n3 B8.n1 152.298
R4220 B8.n6 B8.t8 109.215
R4221 B8.n5 B8.t1 102.659
R4222 B8.n7 B8.n5 47.4474
R4223 B8.n9 B8.n3 19.8357
R4224 B8 B8.n9 15.6269
R4225 B8.n9 B8.n8 1.54462
R4226 A3.n1 A3.t8 373.283
R4227 A3.n0 A3.t9 347.577
R4228 A3.n9 A3.t7 334.723
R4229 A3.n3 A3.t11 323.476
R4230 A3.n3 A3.t0 217.436
R4231 A3.n5 A3.t5 212.081
R4232 A3.n6 A3.t3 212.081
R4233 A3.n9 A3.t1 206.19
R4234 A3.n0 A3.t6 193.337
R4235 A3.n8 A3.n7 174.552
R4236 A3.n4 A3.n3 169.833
R4237 A3.n1 A3.t10 167.63
R4238 A3.n2 A3.n0 166.843
R4239 A3.n2 A3.n1 166.421
R4240 A3.n10 A3.n9 152
R4241 A3.n5 A3.t4 139.78
R4242 A3.n6 A3.t2 139.78
R4243 A3.n7 A3.n6 37.246
R4244 A3.n7 A3.n5 24.1005
R4245 A3.n10 A3.n8 17.5294
R4246 A3.n4 A3.n2 1.55989
R4247 A3 A3.n10 0.914786
R4248 A3.n8 A3.n4 0.112749
R4249 B15.n9 B15.t2 384.529
R4250 B15.n3 B15.t11 373.283
R4251 B15.n5 B15.t1 351.861
R4252 B15.n4 B15.t7 297.233
R4253 B15.n2 B15.n1 257.209
R4254 B15.n0 B15.t4 241.536
R4255 B15.n1 B15.t10 241.536
R4256 B15.n6 B15.n5 214.362
R4257 B15.n0 B15.t3 169.237
R4258 B15.n1 B15.t9 169.237
R4259 B15.n7 B15.n3 167.825
R4260 B15.n3 B15.t8 167.63
R4261 B15.n7 B15.n6 163.79
R4262 B15.n9 B15.t0 156.382
R4263 B15.n2 B15.n0 153.97
R4264 B15.n10 B15.n9 152
R4265 B15.n5 B15.t6 109.215
R4266 B15.n4 B15.t5 102.659
R4267 B15.n6 B15.n4 47.4474
R4268 B15.n8 B15.n2 20.0296
R4269 B15.n10 B15.n8 16.0683
R4270 B15.n8 B15.n7 1.54462
R4271 B15 B15.n10 0.294753
R4272 A0.n1 A0.t9 373.283
R4273 A0.n0 A0.t6 347.577
R4274 A0.n9 A0.t11 334.723
R4275 A0.n3 A0.t1 323.476
R4276 A0.n3 A0.t2 217.436
R4277 A0.n5 A0.t7 212.081
R4278 A0.n6 A0.t3 212.081
R4279 A0.n9 A0.t0 206.19
R4280 A0.n0 A0.t4 193.337
R4281 A0.n8 A0.n7 171.9
R4282 A0.n4 A0.n3 169.833
R4283 A0.n1 A0.t8 167.63
R4284 A0.n2 A0.n0 166.843
R4285 A0.n2 A0.n1 166.421
R4286 A0.n10 A0.n9 152
R4287 A0.n5 A0.t5 139.78
R4288 A0.n6 A0.t10 139.78
R4289 A0.n7 A0.n6 37.246
R4290 A0.n7 A0.n5 24.1005
R4291 A0.n10 A0.n8 17.5294
R4292 A0 A0.n10 1.82907
R4293 A0.n4 A0.n2 1.55989
R4294 A0.n8 A0.n4 0.112749
R4295 B12.n0 B12.t2 384.529
R4296 B12.n4 B12.t6 373.283
R4297 B12.n6 B12.t8 351.861
R4298 B12.n5 B12.t10 297.233
R4299 B12.n3 B12.n2 263.558
R4300 B12.n1 B12.t0 241.536
R4301 B12.n2 B12.t1 241.536
R4302 B12.n7 B12.n6 214.362
R4303 B12.n1 B12.t9 169.237
R4304 B12.n2 B12.t11 169.237
R4305 B12.n8 B12.n4 167.825
R4306 B12.n4 B12.t5 167.63
R4307 B12.n8 B12.n7 163.79
R4308 B12.n0 B12.t4 156.382
R4309 B12 B12.n0 154.649
R4310 B12.n3 B12.n1 152.298
R4311 B12.n6 B12.t3 109.215
R4312 B12.n5 B12.t7 102.659
R4313 B12.n7 B12.n5 47.4474
R4314 B12.n9 B12.n3 19.8357
R4315 B12 B12.n9 13.42
R4316 B12.n9 B12.n8 1.54462
R4317 B5.n9 B5.t1 384.529
R4318 B5.n0 B5.t0 373.283
R4319 B5.n2 B5.t2 351.861
R4320 B5.n1 B5.t9 297.233
R4321 B5.n7 B5.n5 257.209
R4322 B5.n6 B5.t6 241.536
R4323 B5.n5 B5.t10 241.536
R4324 B5.n3 B5.n2 214.362
R4325 B5.n6 B5.t3 169.237
R4326 B5.n5 B5.t5 169.237
R4327 B5.n4 B5.n0 167.825
R4328 B5.n0 B5.t7 167.63
R4329 B5.n4 B5.n3 163.79
R4330 B5.n9 B5.t8 156.382
R4331 B5.n7 B5.n6 153.97
R4332 B5.n10 B5.n9 152
R4333 B5.n2 B5.t11 109.215
R4334 B5.n1 B5.t4 102.659
R4335 B5.n3 B5.n1 47.4474
R4336 B5.n8 B5.n7 20.032
R4337 B5.n10 B5.n8 16.0683
R4338 B5.n8 B5.n4 1.54462
R4339 B5 B5.n10 0.736132
R4340 B4.n9 B4.t7 384.529
R4341 B4.n0 B4.t11 373.283
R4342 B4.n2 B4.t6 351.861
R4343 B4.n1 B4.t0 297.233
R4344 B4.n7 B4.n5 263.558
R4345 B4.n6 B4.t2 241.536
R4346 B4.n5 B4.t3 241.536
R4347 B4.n3 B4.n2 214.362
R4348 B4.n6 B4.t9 169.237
R4349 B4.n5 B4.t10 169.237
R4350 B4.n4 B4.n0 167.825
R4351 B4.n0 B4.t5 167.63
R4352 B4.n4 B4.n3 163.79
R4353 B4.n9 B4.t1 156.382
R4354 B4.n7 B4.n6 152.298
R4355 B4 B4.n9 152
R4356 B4.n2 B4.t4 109.215
R4357 B4.n1 B4.t8 102.659
R4358 B4.n3 B4.n1 47.4474
R4359 B4.n8 B4.n7 19.8357
R4360 B4 B4.n8 16.0683
R4361 B4.n8 B4.n4 1.54462
R4362 S15 S15.t1 244.464
R4363 S15 S15.t0 165.133
R4364 A12.n1 A12.t0 373.283
R4365 A12.n0 A12.t7 347.577
R4366 A12.n9 A12.t5 334.723
R4367 A12.n3 A12.t10 323.476
R4368 A12.n3 A12.t11 217.436
R4369 A12.n5 A12.t6 212.081
R4370 A12.n6 A12.t8 212.081
R4371 A12.n9 A12.t9 206.19
R4372 A12.n0 A12.t3 193.337
R4373 A12.n8 A12.n7 171.9
R4374 A12.n4 A12.n3 169.833
R4375 A12.n1 A12.t2 167.63
R4376 A12.n2 A12.n0 166.843
R4377 A12.n2 A12.n1 166.421
R4378 A12.n10 A12.n9 152
R4379 A12.n5 A12.t1 139.78
R4380 A12.n6 A12.t4 139.78
R4381 A12.n7 A12.n5 37.246
R4382 A12.n7 A12.n6 24.1005
R4383 A12.n10 A12.n8 17.5294
R4384 A12 A12.n10 1.82907
R4385 A12.n4 A12.n2 1.55989
R4386 A12.n8 A12.n4 0.112749
R4387 B11.n9 B11.t1 384.529
R4388 B11.n3 B11.t11 373.283
R4389 B11.n5 B11.t0 351.861
R4390 B11.n4 B11.t5 297.233
R4391 B11.n2 B11.n1 257.209
R4392 B11.n0 B11.t8 241.536
R4393 B11.n1 B11.t3 241.536
R4394 B11.n6 B11.n5 214.362
R4395 B11.n0 B11.t4 169.237
R4396 B11.n1 B11.t10 169.237
R4397 B11.n7 B11.n3 167.825
R4398 B11.n3 B11.t2 167.63
R4399 B11.n7 B11.n6 163.79
R4400 B11.n9 B11.t6 156.382
R4401 B11.n2 B11.n0 153.97
R4402 B11.n10 B11.n9 152
R4403 B11.n5 B11.t7 109.215
R4404 B11.n4 B11.t9 102.659
R4405 B11.n6 B11.n4 47.4474
R4406 B11.n8 B11.n2 20.0296
R4407 B11.n10 B11.n8 16.0683
R4408 B11 B11.n10 1.61889
R4409 B11.n8 B11.n7 1.54462
R4410 Cin.n0 Cin.t2 471.289
R4411 Cin.n1 Cin.t1 373.283
R4412 Cin.n4 Cin.n2 357.442
R4413 Cin.n3 Cin.t4 346.022
R4414 Cin.n2 Cin.t0 325.082
R4415 Cin.n2 Cin.t6 215.829
R4416 Cin Cin.n0 212.018
R4417 Cin.n3 Cin.t7 193.337
R4418 Cin.n1 Cin.t5 167.63
R4419 Cin.n4 Cin.n3 152
R4420 Cin Cin.n1 152
R4421 Cin.n0 Cin.t3 148.35
R4422 Cin Cin.n4 86.1712
R4423 B7.n9 B7.t2 384.529
R4424 B7.n0 B7.t1 373.283
R4425 B7.n2 B7.t3 351.861
R4426 B7.n1 B7.t8 297.233
R4427 B7.n7 B7.n5 257.209
R4428 B7.n6 B7.t9 241.536
R4429 B7.n5 B7.t10 241.536
R4430 B7.n3 B7.n2 214.362
R4431 B7.n6 B7.t4 169.237
R4432 B7.n5 B7.t5 169.237
R4433 B7.n4 B7.n0 167.825
R4434 B7.n0 B7.t6 167.63
R4435 B7.n4 B7.n3 163.79
R4436 B7.n9 B7.t7 156.382
R4437 B7.n7 B7.n6 153.97
R4438 B7.n10 B7.n9 152
R4439 B7.n2 B7.t11 109.215
R4440 B7.n1 B7.t0 102.659
R4441 B7.n3 B7.n1 47.4474
R4442 B7.n8 B7.n7 20.032
R4443 B7.n10 B7.n8 16.0683
R4444 B7 B7.n10 1.61889
R4445 B7.n8 B7.n4 1.54462
R4446 A9.n1 A9.t7 373.283
R4447 A9.n0 A9.t1 347.577
R4448 A9.n9 A9.t6 334.723
R4449 A9.n3 A9.t5 323.476
R4450 A9.n3 A9.t9 217.436
R4451 A9.n5 A9.t2 212.081
R4452 A9.n6 A9.t4 212.081
R4453 A9.n9 A9.t0 206.19
R4454 A9.n0 A9.t8 193.337
R4455 A9.n8 A9.n7 174.552
R4456 A9.n4 A9.n3 169.833
R4457 A9.n1 A9.t3 167.63
R4458 A9.n2 A9.n0 166.843
R4459 A9.n2 A9.n1 166.421
R4460 A9.n10 A9.n9 152
R4461 A9.n5 A9.t10 139.78
R4462 A9.n6 A9.t11 139.78
R4463 A9.n7 A9.n5 37.246
R4464 A9.n7 A9.n6 24.1005
R4465 A9.n10 A9.n8 17.5294
R4466 A9.n4 A9.n2 1.55989
R4467 A9 A9.n10 0.457643
R4468 A9.n8 A9.n4 0.112749
R4469 A5.n1 A5.t1 373.283
R4470 A5.n0 A5.t9 347.577
R4471 A5.n9 A5.t5 334.723
R4472 A5.n3 A5.t3 323.476
R4473 A5.n3 A5.t10 217.436
R4474 A5.n5 A5.t7 212.081
R4475 A5.n6 A5.t6 212.081
R4476 A5.n9 A5.t11 206.19
R4477 A5.n0 A5.t4 193.337
R4478 A5.n8 A5.n7 174.552
R4479 A5.n4 A5.n3 169.833
R4480 A5.n1 A5.t8 167.63
R4481 A5.n2 A5.n0 166.843
R4482 A5.n2 A5.n1 166.421
R4483 A5.n10 A5.n9 152
R4484 A5.n5 A5.t2 139.78
R4485 A5.n6 A5.t0 139.78
R4486 A5.n7 A5.n6 37.246
R4487 A5.n7 A5.n5 24.1005
R4488 A5.n10 A5.n8 17.5294
R4489 A5 A5.n10 2.28621
R4490 A5.n4 A5.n2 1.55989
R4491 A5.n8 A5.n4 0.112749
R4492 B1.n9 B1.t5 384.529
R4493 B1.n0 B1.t2 373.283
R4494 B1.n2 B1.t9 351.861
R4495 B1.n1 B1.t6 297.233
R4496 B1.n7 B1.n5 257.209
R4497 B1.n6 B1.t10 241.536
R4498 B1.n5 B1.t4 241.536
R4499 B1.n3 B1.n2 214.362
R4500 B1.n6 B1.t7 169.237
R4501 B1.n5 B1.t1 169.237
R4502 B1.n4 B1.n0 167.825
R4503 B1.n0 B1.t8 167.63
R4504 B1.n4 B1.n3 163.79
R4505 B1.n9 B1.t0 156.382
R4506 B1.n7 B1.n6 153.97
R4507 B1 B1.n9 152.294
R4508 B1.n2 B1.t3 109.215
R4509 B1.n1 B1.t11 102.659
R4510 B1.n3 B1.n1 47.4474
R4511 B1.n8 B1.n7 20.032
R4512 B1 B1.n8 15.7741
R4513 B1.n8 B1.n4 1.54462
R4514 B3.n9 B3.t1 384.529
R4515 B3.n0 B3.t0 373.283
R4516 B3.n2 B3.t2 351.861
R4517 B3.n1 B3.t3 297.233
R4518 B3.n7 B3.n5 257.209
R4519 B3.n6 B3.t5 241.536
R4520 B3.n5 B3.t8 241.536
R4521 B3.n3 B3.n2 214.362
R4522 B3.n6 B3.t4 169.237
R4523 B3.n5 B3.t7 169.237
R4524 B3.n4 B3.n0 167.825
R4525 B3.n0 B3.t6 167.63
R4526 B3.n4 B3.n3 163.79
R4527 B3.n9 B3.t10 156.382
R4528 B3.n7 B3.n6 153.97
R4529 B3.n10 B3.n9 152
R4530 B3.n2 B3.t11 109.215
R4531 B3.n1 B3.t9 102.659
R4532 B3.n3 B3.n1 47.4474
R4533 B3.n8 B3.n7 20.032
R4534 B3.n10 B3.n8 16.0683
R4535 B3.n8 B3.n4 1.54462
R4536 B3 B3.n10 0.294753
R4537 a_3177_n4294.n0 a_3177_n4294.t5 471.289
R4538 a_3177_n4294.n4 a_3177_n4294.t3 373.283
R4539 a_3177_n4294.n3 a_3177_n4294.n1 357.442
R4540 a_3177_n4294.n2 a_3177_n4294.t7 346.022
R4541 a_3177_n4294.n1 a_3177_n4294.t6 325.082
R4542 a_3177_n4294.n7 a_3177_n4294.t0 294.913
R4543 a_3177_n4294.t1 a_3177_n4294.n7 217.999
R4544 a_3177_n4294.n1 a_3177_n4294.t4 215.829
R4545 a_3177_n4294.n2 a_3177_n4294.t8 193.337
R4546 a_3177_n4294.n6 a_3177_n4294.n0 189.391
R4547 a_3177_n4294.n4 a_3177_n4294.t2 167.63
R4548 a_3177_n4294.n3 a_3177_n4294.n2 152
R4549 a_3177_n4294.n5 a_3177_n4294.n4 152
R4550 a_3177_n4294.n0 a_3177_n4294.t9 148.35
R4551 a_3177_n4294.n5 a_3177_n4294.n3 86.1712
R4552 a_3177_n4294.n7 a_3177_n4294.n6 35.6311
R4553 a_3177_n4294.n6 a_3177_n4294.n5 22.6709
C0 a_3946_n1066# B14 3.07e-19
C1 DVDD a_894_n1194# 8.89e-20
C2 a_1557_46# a_1997_46# 0.046215f
C3 a_1201_n574# a_3669_n342# 6.3e-20
C4 a_n131_n574# a_3765_n600# 4.08e-20
C5 a_1557_n1194# a_n131_n1814# 0.002594f
C6 a_636_n1814# a_2908_n600# 0.00211f
C7 a_4204_n3054# a_4363_n2068# 1.97e-19
C8 A15 a_3861_n3080# 1.7e-21
C9 A14 a_5402_174# 0.003407f
C10 a_143_n1036# a_1997_n828# 5.14e-19
C11 DVDD a_5456_412# 0.156886f
C12 a_2273_n254# a_1641_n828# 0.001272f
C13 B3 a_2908_n600# 1.85e-19
C14 DVDD a_2569_n3928# 2.55e-19
C15 B8 a_3861_n3080# 0.059236f
C16 a_3946_174# a_4000_412# 0.004411f
C17 a_3874_20# a_4363_412# 0.12395f
C18 a_147_n254# a_n131_n574# 0.002789f
C19 a_143_n1036# a_n71_n600# 0.001762f
C20 DVDD a_143_n1036# 0.789516f
C21 a_143_n2276# a_1647_n3054# 2.86e-19
C22 a_1997_n3674# a_2273_n2734# 0.001323f
C23 a_3874_n2460# a_4523_n3054# 2.35e-19
C24 a_143_n2276# a_1479_n1494# 6.56e-19
C25 a_636_n574# a_3904_46# 2.15e-20
C26 a_5192_n3674# B10 6.11e-20
C27 B2 a_966_n1194# 6.11e-20
C28 a_3874_n1220# a_4363_n1194# 0.033252f
C29 a_2254_n1194# a_1968_n1814# 1.54e-19
C30 a_798_n1194# a_1557_n1194# 0.031298f
C31 a_3874_n1220# A3 3.62e-21
C32 a_147_n1494# a_n131_n1814# 0.002687f
C33 a_4441_n1814# a_3543_n342# 0.011053f
C34 a_3655_n1516# a_3669_n342# 0.024621f
C35 a_3434_n1546# a_3765_n600# 1.81e-21
C36 a_143_n2276# a_894_n2434# 4.02e-19
C37 A4 a_1261_n3080# 6.77e-21
C38 DVDD a_2569_n1775# 0.108858f
C39 B2 a_2273_n254# 2.25e-20
C40 S15 a_1201_n574# 4.87e-19
C41 a_3434_n4026# a_3904_n3674# 1.54e-19
C42 a_3226_n4062# a_n131_n4294# 5.42e-19
C43 B15 a_4697_n828# 4.23e-20
C44 a_3765_n3080# a_4691_n2734# 0.004527f
C45 a_143_n2276# a_3226_n4062# 0.00255f
C46 a_3669_n2822# a_3904_n3674# 0.023649f
C47 a_4441_n1814# a_4441_n574# 0.002078f
C48 A3 a_n71_n1840# 1.38e-21
C49 a_3322_n1582# a_n131_n574# 1.64e-19
C50 A10 a_4441_n4294# 6.77e-21
C51 B4 a_n131_n1814# 0.015549f
C52 a_5855_n1814# a_3669_n342# 1.83e-19
C53 a_636_n3054# a_n131_n1814# 0.001496f
C54 a_6023_n1814# a_3543_n342# 0.096176f
C55 A10 a_3861_n3080# 2.3e-19
C56 A12 a_3861_n600# 0.025968f
C57 a_1641_n3674# B5 2.95e-21
C58 a_1201_n1814# a_1261_n3080# 4.02e-20
C59 B12 a_5360_n1194# 1.17e-20
C60 A8 a_5456_n2434# 0.047225f
C61 a_3946_n2306# a_3434_n1546# 5.1e-20
C62 a_3874_n2460# a_3655_n1516# 8.78e-19
C63 a_2995_n4294# a_3226_n1582# 0.011655f
C64 A4 a_798_n3674# 2.18e-20
C65 a_636_n574# a_315_n574# 3.68e-19
C66 A12 a_5360_46# 0.114467f
C67 B12 a_5288_412# 3.03e-19
C68 a_798_n2434# A5 0.001236f
C69 A7 a_1968_n4294# 0.00356f
C70 a_1291_n1814# a_636_n1814# 6.24e-19
C71 a_1997_n1194# a_1557_46# 7.6e-20
C72 a_3832_46# a_4000_46# 2.18e-19
C73 a_2995_n4294# a_4000_n2434# 0.005807f
C74 a_3946_n2306# a_4363_n2434# 0.06777f
C75 a_2254_n2434# A9 9.68e-20
C76 a_1291_n1814# B3 0.056553f
C77 A1 a_1261_n600# 0.076981f
C78 a_798_n1194# B4 1.22e-20
C79 A0 A1 0.019542f
C80 B1 a_n71_n600# 3.52e-21
C81 DVDD B1 0.565768f
C82 B0 Cin 0.669312f
C83 A11 a_4000_n3674# 0.046632f
C84 a_3322_n1582# a_3434_n1546# 0.14976f
C85 a_1557_n2434# A3 2.88e-19
C86 a_1997_n2434# a_1557_n1194# 6.4e-20
C87 B5 a_2422_n2434# 6.11e-20
C88 A3 a_1997_46# 6.84e-21
C89 a_n41_n1814# a_n71_n1840# 0.025037f
C90 a_1557_n2434# B9 2.32e-20
C91 a_1479_n1494# a_1968_n1814# 3.05e-19
C92 A9 a_3904_n3674# 2.18e-20
C93 DVDD a_4523_n4294# 0.008551f
C94 A0 a_185_n1194# 1.17e-19
C95 a_4000_n828# a_4363_n828# 0.009846f
C96 a_1641_n828# a_1997_n828# 0.009846f
C97 a_2790_n3928# a_1968_n4294# 3.89e-19
C98 A6 a_n131_n1814# 8.62e-20
C99 a_3434_n4026# a_2273_n2734# 1.42e-19
C100 a_185_n3674# A4 1.17e-19
C101 a_6153_n3674# a_3543_n2822# 1.33e-19
C102 A7 a_1641_n3674# 0.051667f
C103 a_541_412# a_894_412# 2.18e-19
C104 a_3669_n2822# a_2273_n2734# 7.77e-20
C105 DVDD a_1641_n828# 0.160791f
C106 a_5819_n2068# a_5402_n2306# 0.030161f
C107 a_4691_n1814# a_3322_n1582# 1.57e-19
C108 DVDD a_1557_n3674# 0.379168f
C109 A12 a_4204_n574# 0.002173f
C110 a_5288_n828# a_3543_n342# 3.32e-20
C111 a_1557_n1194# a_1201_n1814# 0.044539f
C112 a_5360_n1194# a_2908_n600# 2.38e-20
C113 a_5402_174# a_5819_412# 0.030161f
C114 a_798_n2434# B6 1.22e-20
C115 a_101_n1194# a_1557_n1194# 0.003292f
C116 a_101_n2434# a_n71_n3080# 0.003994f
C117 a_143_n1036# a_185_46# 1.55e-21
C118 a_1291_n4294# a_143_n3516# 1.59e-20
C119 a_3861_n600# a_3904_n2434# 3.7e-21
C120 a_3543_n342# a_4697_n2068# 3.89e-20
C121 a_2995_n4294# a_3627_n2734# 0.001103f
C122 a_3946_n2306# a_3711_n2734# 3.34e-19
C123 A6 a_11_n3674# 4.78e-19
C124 a_636_n1814# B3 1.25417f
C125 B7 a_2350_n3308# 2.91e-19
C126 a_798_n2434# a_143_n3516# 0.002098f
C127 a_4441_n4294# a_2995_n4294# 7.93e-19
C128 A15 a_4363_n1194# 0.051667f
C129 a_101_46# a_1201_n574# 0.003561f
C130 a_4204_n3054# a_5456_n2434# 7.7e-21
C131 A3 A15 0.006192f
C132 a_5402_n2306# a_3765_n3080# 0.003561f
C133 a_3874_n2460# a_5773_n3054# 0.063303f
C134 a_3946_n2306# a_4441_n3054# 0.002379f
C135 a_2995_n4294# a_3861_n3080# 0.008798f
C136 a_n131_n574# a_1261_n1840# 9.27e-21
C137 B7 a_3904_n3674# 1.77e-20
C138 a_5360_n1194# a_5192_n1194# 0.00792f
C139 a_1997_n2434# a_636_n3054# 0.045338f
C140 a_1641_n2434# a_1557_n2434# 0.06777f
C141 B2 a_n71_n600# 0.001373f
C142 DVDD B2 0.822861f
C143 B1 B13 0.001479f
C144 A0 A2 0.009427f
C145 A15 B9 0.00374f
C146 B15 A9 0.007762f
C147 A4 B4 1.27934f
C148 a_101_n2434# a_541_n3308# 4.9e-19
C149 a_636_n3054# A4 0.021138f
C150 a_3946_n1066# a_3434_n1546# 0.116264f
C151 a_3874_n1220# a_3655_n1516# 9.72e-19
C152 a_1201_n1814# a_1647_n574# 1.02e-20
C153 a_1647_n4294# a_2995_n4294# 1.68e-19
C154 a_636_n1814# a_1291_n574# 1.21e-19
C155 a_3711_n254# a_3669_n342# 0.001239f
C156 a_3946_n2306# a_4000_n2068# 0.004411f
C157 a_3711_n2734# a_1201_n3054# 9.58e-21
C158 a_3627_n2734# a_1201_n4294# 2.72e-21
C159 a_3874_n2460# a_4363_n2068# 0.12395f
C160 a_2543_n2734# a_n131_n4294# 2.77e-20
C161 a_3627_n254# a_3765_n600# 3.31e-19
C162 a_2995_n4294# a_3904_n2434# 0.052026f
C163 B9 B8 0.003904f
C164 a_143_n2276# a_2543_n2734# 7.9e-19
C165 DVDD a_2422_n2068# 6.64e-19
C166 DVDD a_3736_n3308# 6.64e-19
C167 B8 a_5192_n2434# 6.11e-20
C168 B4 a_185_n3308# 5.74e-19
C169 B3 a_1291_n574# 0.001447f
C170 a_3874_n3700# a_4363_n3308# 0.12395f
C171 a_3946_n3546# a_4000_n3308# 0.004914f
C172 A8 a_5773_n1814# 0.001911f
C173 a_3861_n3080# a_1201_n4294# 6.1e-20
C174 a_3765_n3080# a_n131_n4294# 3.23e-20
C175 a_n131_n574# a_2254_46# 3.5e-19
C176 a_143_n2276# a_3765_n3080# 1.95e-20
C177 a_636_n3054# a_1201_n1814# 6.57e-20
C178 DVDD a_315_n3054# 0.006628f
C179 B7 a_1261_n4320# 0.2191f
C180 a_101_n1194# B4 3.81e-20
C181 a_1997_n1194# A3 0.046632f
C182 DVDD a_4363_n3308# 0.160791f
C183 a_636_n1814# a_101_n2434# 8.25e-20
C184 a_3874_n1220# a_5855_n1814# 8e-20
C185 A12 a_5402_n1066# 6.66e-20
C186 B12 a_5773_n574# 0.226175f
C187 a_2273_n254# a_2422_46# 2.27e-20
C188 B11 a_3736_n3674# 6.11e-20
C189 a_3226_n4062# a_3685_n4255# 6.64e-19
C190 a_1647_n4294# a_1201_n4294# 0.002223f
C191 a_1291_n4294# a_n131_n4294# 0.017157f
C192 DVDD a_1641_46# 0.001386f
C193 B0 a_966_46# 6.11e-20
C194 Cin a_894_46# 2.5e-19
C195 A14 a_5456_46# 2.43e-21
C196 A10 a_6153_n3308# 5.12e-20
C197 A7 a_3543_n2822# 1.12e-19
C198 A6 A4 0.009427f
C199 a_798_n2434# a_143_n2276# 0.098896f
C200 Cin a_2908_n600# 0.076749f
C201 a_5855_n3054# a_4204_n3054# 8.43e-19
C202 B7 a_2273_n2734# 0.040998f
C203 a_2569_n4255# a_1557_n3674# 4.55e-19
C204 a_4441_n1814# a_4691_n1494# 0.007234f
C205 a_3226_n1582# a_3685_n1775# 6.64e-19
C206 a_3832_n1194# a_4000_n1194# 2.18e-19
C207 DVDD a_1968_n4294# 0.301739f
C208 A6 a_185_n3308# 0.011602f
C209 a_3832_n3674# a_3322_n4062# 4.97e-19
C210 a_3322_n1582# a_3627_n254# 7.04e-19
C211 a_2569_n3928# a_3434_n4026# 3.16e-20
C212 a_2908_n600# a_3669_n342# 0.038268f
C213 a_n131_n1814# a_3765_n600# 3.23e-20
C214 a_147_n2734# a_n131_n1814# 2.42e-19
C215 a_2497_n1775# a_2569_n1775# 6.64e-19
C216 a_5819_n3674# a_5402_n3546# 0.067562f
C217 a_11_n3308# a_143_n3516# 1.23e-20
C218 a_143_n2276# a_2459_n254# 6.17e-20
C219 a_1641_n1194# a_143_n1036# 9.15e-19
C220 Cin a_3874_20# 1.28e-20
C221 A1 a_1557_46# 0.792469f
C222 A8 a_4204_n3054# 0.002173f
C223 a_1997_n3674# a_1557_n3674# 0.046215f
C224 DVDD a_2459_n2734# 1.88e-19
C225 a_147_n254# a_n131_n1814# 6.93e-20
C226 B1 a_2422_412# 3.18e-19
C227 a_636_n574# a_1261_n600# 0.01589f
C228 A0 a_636_n574# 0.021138f
C229 B0 a_101_46# 0.181244f
C230 a_3543_n342# a_5288_n1194# 1.41e-19
C231 DVDD a_1641_n3674# 0.001386f
C232 B14 a_5402_n2306# 5.99e-19
C233 B0 a_n71_n1840# 8.21e-21
C234 a_1467_n2434# A5 5.03e-19
C235 a_3874_n1220# a_4363_n2068# 1.77e-21
C236 a_3946_n1066# a_4000_n2068# 4.48e-19
C237 a_3874_20# a_3669_n342# 7.1e-20
C238 a_3874_n2460# a_2908_n600# 1.34e-20
C239 B2 a_185_46# 8.1e-22
C240 A2 a_541_46# 2.43e-21
C241 A11 A10 0.019542f
C242 a_541_n2068# a_143_n1036# 6.58e-21
C243 B9 a_3861_n600# 1.71e-21
C244 A8 a_5360_n1194# 1.29e-20
C245 a_3543_n342# a_5819_n2434# 0.001123f
C246 S15 a_2908_n600# 0.054669f
C247 A15 a_3655_n1516# 0.002825f
C248 B5 a_2254_n1194# 8.43e-21
C249 A8 a_5192_n2068# 1.05e-19
C250 DVDD a_185_n828# 0.165024f
C251 a_5192_n1194# a_5456_n1194# 8.12e-20
C252 a_3874_20# a_5773_n574# 0.063303f
C253 a_3322_n1582# a_n131_n1814# 4.14e-19
C254 a_4204_n574# a_4000_412# 1.25e-20
C255 a_2995_n4294# a_4363_n1194# 9.13e-19
C256 DVDD a_4363_n828# 0.160791f
C257 B11 a_4204_n3054# 0.020606f
C258 a_n131_n1814# a_1201_n3054# 6.14e-21
C259 a_315_n574# a_143_n1036# 8.43e-19
C260 a_2995_n4294# B9 0.140464f
C261 a_143_n2276# a_2422_n828# 4.67e-20
C262 a_11_n3308# a_n131_n4294# 9e-21
C263 a_3946_174# a_3711_n254# 3.34e-19
C264 B12 a_3946_174# 3.07e-19
C265 a_4204_n574# a_4363_n1194# 9.15e-19
C266 a_2995_n4294# a_5192_n2434# 5.28e-19
C267 B1 a_1641_n1194# 2.95e-21
C268 a_1968_n4294# a_2569_n4255# 0.190276f
C269 DVDD a_3589_n1448# 2.55e-19
C270 DVDD a_5360_n2434# 0.234243f
C271 a_3589_n3928# a_2995_n4294# 0.004112f
C272 B1 a_3904_46# 1.77e-20
C273 a_1467_n2434# a_143_n3516# 9.38e-21
C274 a_3669_n2822# a_4523_n4294# 0.002223f
C275 a_3543_n2822# a_4691_n4294# 0.017157f
C276 a_1467_n2068# a_1557_n2434# 0.006823f
C277 a_1641_n2068# a_636_n3054# 0.12395f
C278 A4 a_147_n2734# 0.001052f
C279 A7 a_3946_n3546# 2.18e-20
C280 a_3322_n1582# a_3832_46# 6.08e-20
C281 a_6023_n3054# a_3543_n342# 5.44e-19
C282 Cin a_636_n1814# 5.66e-19
C283 a_3669_n2822# a_1557_n3674# 9.92e-21
C284 a_3543_n2822# a_3874_n3700# 0.044377f
C285 B5 a_1647_n3054# 0.007771f
C286 Cin B3 2.79e-19
C287 DVDD A14 0.495937f
C288 A1 A3 0.002462f
C289 DVDD a_3543_n2822# 0.911806f
C290 a_1201_n574# a_3861_n600# 4.08e-20
C291 a_1201_n1814# a_3765_n600# 6.3e-20
C292 a_143_n2276# a_3368_n3928# 3.11e-19
C293 A11 a_2995_n4294# 0.009643f
C294 a_3946_n1066# a_n131_n1814# 1.19e-20
C295 a_1557_n1194# a_3543_n342# 1.19e-20
C296 a_3874_n1220# a_2908_n600# 0.069174f
C297 a_636_n1814# a_3669_n342# 1.36e-21
C298 a_1641_n2434# a_2995_n4294# 4.99e-19
C299 a_1557_46# a_1467_46# 0.006958f
C300 B12 a_6023_n1494# 2.47e-20
C301 B13 a_4363_n828# 9.06e-20
C302 a_4204_n3054# a_5192_n2068# 2.91e-20
C303 a_143_n1036# a_2350_n828# 1.19e-20
C304 a_101_46# a_894_46# 3.78e-19
C305 a_2273_n254# a_2254_n1194# 0.023518f
C306 B3 a_3669_n342# 1.03e-20
C307 DVDD a_n41_n4294# 0.265726f
C308 a_n71_n3080# a_n131_n3054# 0.211818f
C309 a_3946_174# a_2908_n600# 3.32e-20
C310 B8 a_5773_n3054# 0.226175f
C311 A13 a_3736_46# 7.66e-19
C312 a_185_n2434# B4 0.021045f
C313 a_3874_n2460# a_5855_n3054# 3.68e-19
C314 a_2995_n4294# a_4523_n3054# 6.46e-19
C315 A15 a_4363_n2068# 1.58e-21
C316 a_143_n2276# a_2790_n1448# 7.89e-19
C317 Cin a_1291_n574# 6.63e-20
C318 a_5288_n828# a_5456_n828# 2.18e-19
C319 a_5456_n3674# B10 0.005557f
C320 a_3543_n342# a_6153_n1194# 1.33e-19
C321 a_n131_n1814# a_1261_n1840# 0.011053f
C322 a_5402_n1066# a_4363_n1194# 1.11e-20
C323 a_3946_n1066# a_4697_n1194# 0.006958f
C324 a_3874_n1220# a_5192_n1194# 3.15e-19
C325 a_1641_n3674# a_1997_n3674# 0.008475f
C326 A12 a_5192_412# 1.05e-19
C327 A11 a_1201_n4294# 7.21e-20
C328 B14 a_6023_n574# 3.35e-19
C329 a_5773_n1814# a_3669_n342# 3.93e-19
C330 a_3655_n1516# a_3861_n600# 5.6e-20
C331 a_4441_n1814# a_3765_n600# 7.34e-21
C332 DVDD a_185_n2068# 0.164242f
C333 a_3874_n1220# a_3874_20# 8.69e-20
C334 a_2350_n3674# a_2995_n4294# 1.05e-19
C335 a_143_n2276# a_1467_n2434# 1.09e-20
C336 A4 a_1201_n3054# 4.94e-20
C337 a_3736_n3308# a_3669_n2822# 1.98e-19
C338 Cin a_2783_n1775# 1.1e-19
C339 A7 a_1647_n3054# 3.39e-19
C340 a_3874_20# a_3946_174# 0.287408f
C341 A8 a_5456_n1194# 2.43e-21
C342 a_636_n574# a_1557_46# 0.287408f
C343 a_3861_n3080# a_6023_n2734# 0.002789f
C344 a_101_n3674# a_n71_n3080# 5.92e-19
C345 a_4441_n3054# a_4691_n2734# 0.007234f
C346 a_3669_n2822# a_4363_n3308# 3.93e-19
C347 A3 a_2315_n1775# 0.002825f
C348 a_3861_n3080# a_3904_n3674# 3.29e-19
C349 a_3322_n1582# a_1201_n1814# 6.64e-20
C350 a_5773_n1814# a_5773_n574# 0.001197f
C351 a_2254_n2434# a_3904_n2434# 0.004465f
C352 a_3874_n2460# A8 0.021138f
C353 a_n131_n1814# a_3368_n1775# 3.15e-20
C354 A2 A3 0.019542f
C355 a_5402_n2306# B10 1.3e-19
C356 A10 a_5773_n3054# 0.001913f
C357 B11 a_4697_n3674# 6.45e-19
C358 A6 a_185_n2434# 4.33e-21
C359 a_1201_n1814# a_1201_n3054# 3.32e-21
C360 a_3946_n2306# a_4441_n1814# 1.81e-19
C361 A8 a_6153_n2434# 4.78e-19
C362 a_2995_n4294# a_3655_n1516# 0.006008f
C363 a_2350_n3674# a_1201_n4294# 6.23e-20
C364 a_143_n2276# a_n131_n574# 0.002272f
C365 B12 a_5819_n828# 5.74e-19
C366 a_541_n3308# a_894_n3308# 2.18e-19
C367 a_3874_20# a_4523_n574# 2.35e-19
C368 A13 a_4363_46# 0.051667f
C369 B7 a_1557_n3674# 0.175017f
C370 a_101_n3674# a_541_n3308# 0.004108f
C371 a_1968_n4294# a_3434_n4026# 0.001915f
C372 a_5402_n2306# a_4363_n2434# 1.11e-20
C373 a_2569_n4255# a_3543_n2822# 5.42e-19
C374 A1 a_1201_n574# 0.081374f
C375 a_3322_n1582# a_4441_n1814# 6.23e-19
C376 a_n71_n3080# a_n71_n1840# 0.001197f
C377 a_3874_n3700# a_5855_n4294# 8e-20
C378 a_2790_n1448# a_1968_n1814# 3.89e-19
C379 DVDD a_5855_n4294# 0.008765f
C380 A9 a_4363_n3308# 1.58e-21
C381 a_1997_n828# a_2254_n1194# 0.02283f
C382 a_1557_46# a_2350_46# 3.53e-19
C383 a_1647_n4294# a_1261_n4320# 0.006406f
C384 a_3177_n1814# a_3226_n1582# 0.077637f
C385 a_143_n2276# a_3434_n1546# 7.28e-19
C386 A2 a_n41_n1814# 0.007489f
C387 a_3874_n3700# a_3946_n3546# 0.287345f
C388 B14 a_5402_174# 1.3e-19
C389 a_3861_n3080# a_2273_n2734# 1.64e-19
C390 DVDD a_2254_n1194# 0.248898f
C391 DVDD a_5819_412# 0.163585f
C392 DVDD a_3946_n3546# 0.379168f
C393 A15 a_2908_n600# 0.118034f
C394 A12 a_6023_n254# 0.001052f
C395 a_3874_20# a_4697_412# 7.45e-20
C396 a_3946_174# a_4363_412# 0.030161f
C397 a_3946_n1066# a_1201_n1814# 9.92e-21
C398 a_3736_n3674# a_4000_n3674# 8.12e-20
C399 a_5456_n828# a_3543_n342# 5.55e-19
C400 A0 a_143_n1036# 0.002173f
C401 a_143_n1036# a_1261_n600# 0.073551f
C402 a_1479_n254# a_n131_n574# 9.28e-20
C403 a_636_n1814# a_3874_n1220# 1.96e-19
C404 B15 a_3904_n2434# 8.78e-21
C405 a_5360_n3674# a_3874_n3700# 0.012687f
C406 a_1647_n4294# a_2273_n2734# 3.9e-20
C407 a_101_n2434# a_n131_n3054# 0.004436f
C408 a_636_n3054# a_1261_n3080# 0.01589f
C409 a_3543_n342# a_5288_n2068# 2.73e-20
C410 a_5402_174# a_4363_46# 1.11e-20
C411 a_3874_n2460# a_4204_n3054# 0.102258f
C412 a_2995_n4294# a_3795_n2734# 0.001418f
C413 a_3946_n2306# a_3322_n4062# 0.008526f
C414 a_3874_n1220# B3 4.99e-21
C415 DVDD a_5360_n3674# 0.234243f
C416 a_966_n2068# a_143_n3516# 2.91e-20
C417 a_3874_n1220# A8 4.8e-19
C418 a_5402_n2306# a_4441_n3054# 0.005909f
C419 a_2995_n4294# a_5773_n3054# 1.52e-19
C420 a_1201_n574# a_2315_n1775# 2.4e-19
C421 a_n131_n574# a_1968_n1814# 5.85e-21
C422 a_1201_n1814# a_1261_n1840# 0.188936f
C423 a_5360_n2434# a_5456_n2068# 0.02283f
C424 a_5360_n1194# a_5456_n1194# 0.023012f
C425 a_101_n1194# a_1261_n1840# 0.005934f
C426 a_636_n1814# a_n71_n1840# 0.062036f
C427 a_1997_n2068# a_n131_n1814# 0.001046f
C428 a_3322_n1582# a_3322_n4062# 6.99e-20
C429 B4 a_798_n3674# 1.17e-20
C430 a_3946_n1066# a_4441_n1814# 0.003171f
C431 a_3874_n1220# a_5773_n1814# 0.062036f
C432 B3 a_n71_n1840# 3.52e-21
C433 a_3832_n3308# a_3946_n3546# 4.35e-21
C434 A5 a_n131_n1814# 8.47e-19
C435 a_3795_n254# a_3765_n600# 0.006083f
C436 a_3946_n2306# a_4697_n2068# 0.006823f
C437 a_3322_n4062# a_1201_n3054# 3.67e-20
C438 a_2995_n4294# a_4363_n2068# 0.016491f
C439 B12 a_3861_n600# 0.059236f
C440 DVDD a_3832_n2068# 4.94e-19
C441 a_101_n2434# a_101_n3674# 0.007891f
C442 B8 a_5456_n2434# 0.005557f
C443 a_3946_n3546# a_4697_n3308# 0.006823f
C444 B12 a_5360_46# 0.078639f
C445 A12 a_5456_412# 0.011819f
C446 a_3322_n1582# a_5288_n828# 1.6e-20
C447 a_1201_n1814# a_2254_46# 3.97e-19
C448 a_3226_n1582# a_2569_n1775# 0.011879f
C449 a_798_n2434# B5 2.55e-19
C450 a_3434_n1546# a_1968_n1814# 0.001915f
C451 a_5456_n2068# A14 3.08e-21
C452 B7 a_1968_n4294# 0.002893f
C453 DVDD a_1647_n3054# 0.005567f
C454 a_2422_n1194# A3 7.66e-19
C455 DVDD a_5192_n3308# 6.64e-19
C456 DVDD a_1479_n1494# 4.62e-19
C457 a_1557_n1194# a_636_n3054# 0.002572f
C458 DVDD a_185_412# 0.165024f
C459 a_2254_n2434# B9 1.77e-20
C460 B11 a_4000_n3674# 0.005557f
C461 B0 A1 1.74e-19
C462 B1 a_1261_n600# 0.214186f
C463 A0 B1 2.69e-19
C464 a_1557_n2434# B3 3.5e-19
C465 a_4441_n1814# a_4691_n574# 9.75e-20
C466 A6 a_798_n3674# 0.114467f
C467 a_966_n2068# a_143_n2276# 5.05e-19
C468 a_101_n2434# a_n71_n1840# 5.92e-19
C469 a_3434_n4026# a_3543_n2822# 0.031799f
C470 a_636_n4294# a_3322_n4062# 7.5e-21
C471 B6 a_n131_n1814# 2.66e-19
C472 a_3543_n2822# a_3669_n2822# 1.11131f
C473 a_5773_n1814# a_6023_n1494# 0.007234f
C474 DVDD a_3226_n4062# 0.105346f
C475 B7 a_1641_n3674# 0.019568f
C476 a_541_412# a_966_412# 1.31e-19
C477 a_798_46# a_894_412# 0.004869f
C478 A7 a_1291_n4294# 0.007493f
C479 A10 a_5456_n2434# 2.43e-21
C480 a_4000_n3674# a_4204_n3054# 4.76e-20
C481 a_3322_n1582# a_3795_n254# 0.010797f
C482 B12 a_4204_n574# 0.002602f
C483 a_2908_n600# a_3861_n600# 5.58e-19
C484 a_3543_n342# a_3765_n600# 6.83e-19
C485 a_143_n3516# a_n131_n1814# 1.24e-19
C486 a_5360_n2434# A9 0.001236f
C487 a_5402_174# a_6153_412# 0.006823f
C488 a_143_n1036# a_541_46# 7.7e-21
C489 B8 a_5855_n3054# 0.007771f
C490 B6 a_11_n3674# 3.15e-19
C491 A6 a_185_n3674# 0.050725f
C492 a_636_n1814# A15 3.62e-21
C493 a_636_n3054# B4 0.014043f
C494 a_4441_n574# a_3765_n600# 0.243071f
C495 a_101_n2434# a_1557_n2434# 0.003292f
C496 B15 a_4363_n1194# 0.019568f
C497 a_636_n574# a_1201_n574# 0.104793f
C498 a_3874_n1220# a_5360_n1194# 0.012687f
C499 a_3543_n342# a_5819_n1194# 0.001149f
C500 A3 B15 2.72e-20
C501 B3 A15 2.72e-20
C502 A11 a_3904_n3674# 0.114346f
C503 a_1997_n2434# A5 0.046632f
C504 a_3874_20# a_3861_n600# 0.289331f
C505 B0 A2 1.68e-19
C506 Cin S15 0.016205f
C507 A0 B2 1.48e-19
C508 a_3946_n2306# a_3543_n342# 0.001955f
C509 a_2995_n4294# a_2908_n600# 0.003679f
C510 a_3874_n2460# a_3669_n342# 6.57e-20
C511 A4 A5 0.019542f
C512 B15 B9 0.004788f
C513 A9 a_3543_n2822# 1.84e-20
C514 a_3874_20# a_5360_46# 0.012687f
C515 A8 B8 1.27934f
C516 a_541_n2434# a_894_n2434# 2.18e-19
C517 S15 a_3669_n342# 6.37e-19
C518 A15 a_5773_n1814# 1.38e-21
C519 a_2350_n1194# a_1201_n1814# 6.23e-20
C520 a_541_n2068# a_185_n2068# 0.009846f
C521 a_2254_n3674# a_2422_n3674# 0.00792f
C522 a_1997_n1194# a_636_n1814# 0.045338f
C523 a_1557_46# a_143_n1036# 0.057421f
C524 a_4204_n574# a_2908_n600# 2.11e-19
C525 a_3322_n1582# a_3543_n342# 0.034838f
C526 B8 a_5773_n1814# 0.001358f
C527 A5 a_1201_n1814# 1.38e-19
C528 a_1997_n1194# B3 0.005557f
C529 DVDD a_5192_n828# 6.64e-19
C530 A6 B4 1.68e-19
C531 A6 a_636_n3054# 4.45e-19
C532 a_n131_n1814# a_n131_n4294# 3.71e-20
C533 a_2995_n4294# a_3874_20# 1.69e-20
C534 B12 a_5402_n1066# 6.9e-19
C535 a_2459_n254# a_2273_n254# 7.42e-19
C536 a_143_n2276# a_n131_n1814# 0.571837f
C537 a_n71_n4320# A4 2.8e-21
C538 a_3322_n1582# a_4441_n574# 6.57e-19
C539 Cin a_966_46# 2.76e-19
C540 a_5360_n2434# a_5402_n3546# 9.75e-22
C541 A14 a_5819_46# 4.33e-21
C542 a_5402_n2306# a_5288_n2434# 3.78e-19
C543 a_2995_n4294# a_5456_n2434# 0.045338f
C544 a_4204_n574# a_5192_n1194# 1.32e-19
C545 B6 A4 1.48e-19
C546 B7 a_3543_n2822# 1.25e-20
C547 a_2569_n4255# a_3226_n4062# 0.011879f
C548 DVDD a_5819_n2068# 0.162119f
C549 a_2783_n4255# a_2995_n4294# 3.93e-19
C550 A1 a_2908_n600# 1.93e-19
C551 a_3874_20# a_4204_n574# 0.102258f
C552 a_4441_n4294# a_4523_n4294# 0.006406f
C553 a_1997_n2434# a_143_n3516# 7.87e-20
C554 a_3543_n2822# a_6023_n4294# 0.096176f
C555 A10 A8 0.009427f
C556 a_3669_n2822# a_5855_n4294# 1.83e-19
C557 a_11_n3674# a_n131_n4294# 1.33e-19
C558 A4 a_143_n3516# 0.002173f
C559 a_143_n2276# a_798_n1194# 1.34e-20
C560 B6 a_185_n3308# 0.033026f
C561 a_541_n1194# a_n131_n1814# 0.001186f
C562 B12 a_5855_n574# 0.007771f
C563 DVDD a_2543_n2734# 2.46e-19
C564 a_3434_n4026# a_3946_n3546# 0.116264f
C565 a_3655_n3996# a_3874_n3700# 9.72e-19
C566 Cin a_3874_n1220# 1.96e-21
C567 a_3543_n2822# a_5402_n3546# 0.034089f
C568 a_3669_n2822# a_3946_n3546# 0.044539f
C569 a_3765_n3080# a_3874_n3700# 1.04e-19
C570 DVDD a_3655_n3996# 0.1905f
C571 a_185_n3308# a_143_n3516# 0.091015f
C572 a_2497_n4255# a_n131_n4294# 9.8e-19
C573 DVDD a_3765_n3080# 0.180057f
C574 A1 a_3874_20# 2.02e-20
C575 B1 a_1557_46# 0.17279f
C576 Cin a_3946_174# 1.42e-20
C577 a_3946_n1066# a_3543_n342# 0.002594f
C578 B8 a_4204_n3054# 0.002602f
C579 a_3874_n1220# a_3669_n342# 0.105485f
C580 a_2350_n3674# a_2273_n2734# 4.97e-19
C581 Cin a_101_46# 0.221376f
C582 B0 a_636_n574# 0.014043f
C583 a_5456_n3308# a_3543_n2822# 5.55e-19
C584 a_2273_n254# a_2422_n828# 1.91e-19
C585 a_798_n1194# a_541_n1194# 0.023012f
C586 DVDD a_1291_n4294# 0.260214f
C587 a_1261_n3080# a_1201_n3054# 0.243071f
C588 a_1467_n2434# B5 6.45e-19
C589 a_3946_174# a_3669_n342# 0.016609f
C590 A15 a_5360_n1194# 0.001236f
C591 B11 A10 2.69e-19
C592 a_798_n2434# DVDD 0.234243f
C593 a_3946_n1066# a_4441_n574# 1.81e-19
C594 a_6153_n3674# B10 3.15e-19
C595 a_n131_n1814# a_1968_n1814# 0.031799f
C596 B8 a_5360_n1194# 1.22e-20
C597 a_5402_n1066# a_5192_n1194# 3.46e-19
C598 B15 a_3655_n1516# 2.1e-19
C599 B8 a_5192_n2068# 3.18e-19
C600 A3 a_143_n1036# 0.011053f
C601 A0 a_185_n828# 7.78e-19
C602 a_5773_n1814# a_3861_n600# 1.01e-20
C603 DVDD a_541_n828# 0.157566f
C604 a_5402_n1066# a_3874_20# 1.11e-19
C605 A9 a_3946_n3546# 2.88e-19
C606 a_3736_n3674# a_2995_n4294# 2.35e-19
C607 a_3874_n1220# a_3874_n2460# 0.001068f
C608 a_143_n2276# a_1997_n2434# 0.003902f
C609 a_4204_n574# a_4363_412# 1.97e-19
C610 a_3669_n342# a_4523_n574# 1.02e-20
C611 A4 a_n131_n4294# 3.84e-19
C612 a_143_n2276# A4 0.477544f
C613 B5 a_n131_n574# 1.71e-21
C614 a_5402_n1066# a_5456_n2434# 4.36e-20
C615 A10 a_4204_n3054# 0.467991f
C616 DVDD a_2459_n254# 1.88e-19
C617 a_3543_n2822# a_5288_n3308# 3.32e-20
C618 a_101_n3674# a_n131_n3054# 2.05e-19
C619 a_5773_n3054# a_6023_n2734# 0.007234f
C620 Cin a_1997_46# 0.002419f
C621 a_636_n4294# a_1261_n3080# 5.78e-19
C622 a_n41_n574# a_n131_n574# 0.131556f
C623 a_2995_n4294# A8 0.4803f
C624 a_185_n3308# a_n131_n4294# 5.74e-19
C625 a_1557_n1194# a_3322_n1582# 8.35e-21
C626 a_3543_n342# a_3368_n1775# 8.19e-19
C627 a_4441_n574# a_4691_n574# 0.025037f
C628 B4 a_147_n2734# 0.002402f
C629 a_143_n2276# a_185_n3308# 1.77e-21
C630 a_1641_n2068# a_1997_n2068# 0.009846f
C631 a_2995_n4294# a_5773_n1814# 3.57e-20
C632 a_798_n3674# a_966_n3308# 0.007578f
C633 a_143_n2276# a_1201_n1814# 0.133901f
C634 a_143_n2276# a_2422_n3674# 2.14e-20
C635 a_541_n3674# a_101_n2434# 4.36e-20
C636 a_1557_n1194# a_1201_n3054# -5.88e-38
C637 a_143_n2276# a_101_n1194# 0.005011f
C638 a_3874_20# a_5855_n574# 3.68e-19
C639 a_1641_n2068# A5 0.011562f
C640 A4 a_541_n1194# 2.43e-21
C641 a_n41_n1814# a_143_n1036# 1.35e-19
C642 a_1647_n1814# B3 0.007771f
C643 a_101_n3674# a_894_n3308# 4.35e-21
C644 a_636_n4294# a_798_n3674# 0.012687f
C645 a_3226_n4062# a_3434_n4026# 0.190276f
C646 B7 a_3946_n3546# 2.32e-20
C647 a_3226_n4062# a_3669_n2822# 1.29e-20
C648 a_4204_n574# a_5773_n1814# 1.52e-19
C649 A1 a_636_n1814# 0.004204f
C650 a_1261_n3080# a_1261_n1840# 0.002078f
C651 a_n131_n3054# a_n71_n1840# 1.74e-20
C652 a_5288_n3674# a_4204_n3054# 1.28e-19
C653 a_798_n2434# a_541_n2434# 0.023012f
C654 A2 a_n71_n3080# 1.82e-21
C655 B1 A3 0.007762f
C656 A1 B3 0.004004f
C657 Cin A15 1.35e-19
C658 DVDD B14 0.794861f
C659 a_3368_n1448# a_3434_n1546# 3.89e-19
C660 a_1997_n828# a_2422_n828# 1.31e-19
C661 a_2254_n1194# a_2350_n828# 0.004869f
C662 a_143_n2276# a_4441_n1814# 1.37e-19
C663 a_101_n1194# a_541_n1194# 0.044963f
C664 B11 a_2995_n4294# 0.006385f
C665 a_1557_46# a_1641_46# 0.06777f
C666 a_3946_n3546# a_5402_n3546# 0.003292f
C667 a_101_46# a_966_46# 3.46e-19
C668 a_636_n574# a_894_46# 2.34e-19
C669 DVDD a_2422_n828# 6.64e-19
C670 A15 a_3669_n342# 0.077871f
C671 DVDD a_11_n3308# 5.28e-19
C672 A13 a_3832_46# 5.43e-19
C673 B13 a_3736_46# 6.11e-20
C674 DVDD a_4363_46# 0.001386f
C675 a_6153_n828# a_3543_n342# 9e-21
C676 a_636_n574# a_2908_n600# 1.61e-21
C677 a_2273_n254# a_n131_n574# 0.158736f
C678 a_143_n1036# a_1201_n574# 0.068052f
C679 B4 a_1201_n3054# 4.3e-20
C680 a_1557_n1194# a_3946_n1066# 0.001288f
C681 A3 a_1641_n828# 0.011964f
C682 B15 a_4363_n2068# 9.06e-20
C683 a_636_n3054# a_1201_n3054# 0.104793f
C684 a_1557_n2434# a_n131_n3054# 0.060379f
C685 A1 a_1291_n574# 0.007493f
C686 a_5360_n3674# a_5402_n3546# 0.057934f
C687 a_2995_n4294# a_4204_n3054# 0.047933f
C688 a_1997_412# a_2254_46# 0.02283f
C689 a_3226_n1582# a_3543_n2822# 2.63e-20
C690 DVDD a_5819_n3308# 0.162119f
C691 B12 a_5192_412# 3.18e-19
C692 B11 a_1201_n4294# 1.03e-20
C693 Cin a_1997_n1194# 8.49e-20
C694 a_1641_n2068# a_143_n3516# 1.97e-19
C695 a_3874_n1220# a_3946_174# 0.002601f
C696 a_5288_412# a_5360_46# 0.004869f
C697 a_5402_n1066# A8 0.003351f
C698 a_1201_n1814# a_1968_n1814# 0.055436f
C699 a_5360_n3674# a_5456_n3308# 0.02283f
C700 a_5456_n2068# a_5819_n2068# 0.009846f
C701 a_2350_n2068# a_n131_n1814# 2.73e-20
C702 a_101_n1194# a_1968_n1814# 4.58e-20
C703 a_636_n1814# a_2315_n1775# 9.72e-19
C704 a_1557_n1194# a_1261_n1840# 0.003171f
C705 A15 a_3874_n2460# 0.00421f
C706 A2 a_636_n1814# 0.020957f
C707 a_5402_n1066# a_5773_n1814# 0.003994f
C708 a_2995_n4294# a_5360_n1194# 1.34e-20
C709 a_636_n574# a_3874_20# 0.001289f
C710 a_3434_n1546# a_2273_n254# 1.71e-19
C711 DVDD a_3368_n3928# 4.92e-19
C712 B3 a_2315_n1775# 2.1e-19
C713 a_3874_n2460# B8 0.014043f
C714 a_2995_n4294# a_5192_n2068# 4.74e-19
C715 A12 A14 0.009427f
C716 A2 B3 2.69e-19
C717 B2 A3 1.74e-19
C718 a_n131_n1814# a_n41_n3054# 5.44e-19
C719 a_3322_n4062# a_n131_n4294# 3.18e-19
C720 a_143_n2276# a_3322_n4062# 9.49e-19
C721 a_636_n3054# a_636_n4294# 8.69e-20
C722 B6 a_185_n2434# 8.1e-22
C723 B8 a_6153_n2434# 3.15e-19
C724 a_6023_n3974# B8 2.47e-20
C725 a_4204_n574# a_5360_n1194# 0.079554f
C726 a_1557_n1194# a_2254_46# 3.32e-21
C727 DVDD a_2790_n1448# 4.92e-19
C728 B13 a_4363_46# 0.019568f
C729 a_185_n2434# a_143_n3516# 1.55e-21
C730 a_4204_n574# a_5288_412# 3.3e-20
C731 A13 a_4697_46# 5.03e-19
C732 A11 a_1557_n3674# 2.18e-20
C733 B1 a_1201_n574# 0.097286f
C734 a_5456_n3308# a_5192_n3308# 1.31e-19
C735 a_5360_n3674# a_5288_n3308# 0.004869f
C736 A9 a_3832_n2434# 5.43e-19
C737 a_3669_n2822# a_2543_n2734# 2.72e-21
C738 a_3543_n2822# a_3627_n2734# 2.77e-20
C739 a_3434_n4026# a_3655_n3996# 0.153192f
C740 A6 a_966_n3308# 1.05e-19
C741 B9 a_4363_n3308# 9.06e-20
C742 a_1641_n2068# a_143_n2276# 0.013863f
C743 a_1557_46# a_2422_46# 3.12e-19
C744 a_636_n3054# a_1261_n1840# 5.78e-19
C745 a_3655_n3996# a_3669_n2822# 0.024621f
C746 a_3434_n4026# a_3765_n3080# 1.81e-21
C747 a_4441_n4294# a_3543_n2822# 0.011053f
C748 Cin a_3861_n600# 3.22e-20
C749 A3 a_1641_46# 1.4e-21
C750 A10 a_3874_n2460# 4.45e-19
C751 B2 a_n41_n1814# 0.056624f
C752 a_3669_n2822# a_3765_n3080# 0.15552f
C753 a_3543_n2822# a_3861_n3080# 0.001745f
C754 a_101_46# a_1997_46# 5.42e-21
C755 A2 a_101_n2434# 6.58e-20
C756 a_4441_n1814# a_4523_n1814# 0.006406f
C757 A6 a_636_n4294# 0.020957f
C758 DVDD a_6153_412# 5.28e-19
C759 B15 a_2908_n600# 0.07853f
C760 a_3669_n342# a_3861_n600# 0.006573f
C761 B12 a_6023_n254# 0.002402f
C762 A13 a_4441_n1814# 8.18e-21
C763 a_2350_n3674# a_1557_n3674# 2.79e-19
C764 A10 a_6023_n3974# 0.001052f
C765 a_3946_174# a_4697_412# 0.006823f
C766 B0 a_143_n1036# 0.002602f
C767 DVDD a_n131_n574# 1.68401f
C768 a_n71_n600# a_n131_n574# 0.211818f
C769 A5 a_1261_n3080# 0.076981f
C770 a_3874_n1220# A15 0.51166f
C771 A11 a_3736_n3308# 1.05e-19
C772 a_5773_n574# a_3861_n600# 0.211818f
C773 a_5402_n1066# a_5360_n1194# 0.057934f
C774 a_3874_n3700# B10 0.013754f
C775 a_636_n1814# a_636_n574# 8.69e-20
C776 a_3874_n1220# B8 1.83e-19
C777 a_3589_n3928# a_1968_n4294# 3.16e-20
C778 A15 a_3946_174# 3.41e-19
C779 a_143_n2276# a_185_n2434# 0.033252f
C780 A11 a_4363_n3308# 0.011964f
C781 a_4697_n3674# a_2995_n4294# 4.66e-21
C782 DVDD B10 0.784378f
C783 a_2995_n4294# a_3669_n342# 0.014645f
C784 a_5402_n2306# a_3543_n342# 0.015023f
C785 a_3874_n2460# a_3861_n600# 4.68e-22
C786 A9 a_3765_n3080# 0.081374f
C787 A4 a_n41_n3054# 0.007489f
C788 DVDD a_3434_n1546# 0.306924f
C789 a_541_n2068# a_798_n2434# 0.02283f
C790 B5 a_n131_n1814# 7.3e-19
C791 a_3832_n828# a_2908_n600# 0.004979f
C792 a_3874_n3700# a_4363_n2434# 1.55e-21
C793 S15 a_3861_n600# 1.21e-19
C794 a_2254_n2434# a_636_n1814# 1.17e-20
C795 a_1997_n2068# a_1557_n1194# 4.48e-19
C796 a_2783_n4255# a_2273_n2734# 0.006879f
C797 A15 a_4523_n574# 3.39e-19
C798 a_2350_n1194# a_1557_n1194# 2.79e-19
C799 a_4204_n574# a_3669_n342# 0.022242f
C800 a_n41_n574# a_n131_n1814# 4.81e-19
C801 a_3322_n1582# a_3765_n600# 0.202439f
C802 DVDD a_4363_n2434# 0.001386f
C803 a_3904_46# a_3736_46# 0.00792f
C804 B12 a_5456_412# 0.017703f
C805 A12 a_5819_412# 0.011602f
C806 a_2995_n4294# a_5456_n1194# 7.7e-21
C807 a_2254_n2434# B3 8.78e-21
C808 a_636_n574# a_1291_n574# 0.006212f
C809 a_1557_n1194# A5 1.91e-19
C810 a_2422_n1194# B3 6.11e-20
C811 a_3736_n3674# a_3904_n3674# 0.00792f
C812 DVDD a_4691_n1814# 0.259614f
C813 a_3177_n1814# a_2908_n600# 0.001342f
C814 a_143_n2276# a_3543_n342# 0.008482f
C815 a_147_n2734# a_1201_n3054# 2.05e-20
C816 a_143_n3516# a_1261_n3080# 0.073551f
C817 a_1479_n2734# a_n131_n3054# 9.28e-20
C818 a_3874_n2460# a_2995_n4294# 0.237398f
C819 DVDD a_541_412# 0.157566f
C820 A0 a_185_412# 0.011602f
C821 B0 B1 0.003904f
C822 Cin A1 0.047249f
C823 a_4204_n574# a_5773_n574# 0.001762f
C824 a_4691_n254# a_4441_n574# 0.007234f
C825 a_5402_n2306# a_5819_n2434# 0.067562f
C826 a_4204_n574# a_5456_n1194# 0.045338f
C827 a_3322_n4062# a_3685_n4255# 0.005265f
C828 B6 a_798_n3674# 0.078521f
C829 DVDD a_11_n2434# 2.33e-19
C830 A8 a_6023_n2734# 0.001052f
C831 a_143_n3516# a_798_n3674# 0.079554f
C832 a_798_46# a_966_412# 0.007578f
C833 B7 a_1291_n4294# 0.056553f
C834 a_2995_n4294# a_n131_n3054# 0.003746f
C835 a_966_n1194# a_n131_n1814# 1.65e-19
C836 a_5773_n4294# a_3874_n3700# 0.062036f
C837 a_894_n3674# a_798_n3674# 0.005587f
C838 a_4441_n4294# a_3946_n3546# 0.003171f
C839 DVDD a_3711_n2734# 1.88e-19
C840 a_5360_n2434# B9 2.55e-19
C841 a_1997_n2068# a_636_n3054# 0.112124f
C842 a_3861_n3080# a_3946_n3546# 6.4e-19
C843 a_4441_n3054# a_3874_n3700# 5.78e-19
C844 a_1997_n3308# a_1557_n2434# 5.56e-19
C845 a_143_n1036# a_894_46# 1.66e-19
C846 DVDD a_5773_n4294# 0.183389f
C847 a_5360_n2434# a_5192_n2434# 0.00792f
C848 a_541_n3674# a_101_n3674# 0.044963f
C849 DVDD a_4441_n3054# 0.17389f
C850 B6 a_185_n3674# 0.021045f
C851 B4 A5 1.74e-19
C852 a_636_n1814# B15 4.99e-21
C853 a_636_n3054# A5 0.512147f
C854 a_5402_n1066# a_3669_n342# 0.003559f
C855 a_3874_n1220# a_3861_n600# 0.003854f
C856 a_3946_n1066# a_3765_n600# 5.07e-20
C857 a_143_n1036# a_2908_n600# 7.98e-21
C858 a_2273_n254# a_n131_n1814# 0.034838f
C859 a_1997_n2434# a_2350_n2434# 2.18e-19
C860 a_3946_n3546# a_3904_n2434# 3.32e-21
C861 a_6153_n3308# a_3543_n2822# 9e-21
C862 B3 B15 0.001479f
C863 Cin a_2315_n1775# 0.040089f
C864 a_798_n1194# a_966_n1194# 0.00792f
C865 A3 a_1467_n1194# 5.03e-19
C866 a_185_n3674# a_143_n3516# 0.033252f
C867 a_1997_n2434# B5 0.005557f
C868 a_n131_n3054# a_1201_n4294# 0.006573f
C869 B11 a_3904_n3674# 0.077341f
C870 a_143_n2276# a_1261_n3080# 0.002929f
C871 A1 S15 4.85e-21
C872 DVDD a_4000_n2068# 0.154852f
C873 a_3946_174# a_3861_n600# 0.060379f
C874 B0 B2 0.013937f
C875 a_5819_n3674# A8 1.17e-19
C876 A4 B5 2.69e-19
C877 B9 a_3543_n2822# 2.07e-21
C878 a_966_n2068# DVDD 6.64e-19
C879 a_5402_n1066# a_5773_n574# 5.92e-19
C880 a_2908_n600# a_2569_n1775# 7.8e-19
C881 a_3543_n342# a_1968_n1814# 2.79e-19
C882 a_1557_46# a_2254_n1194# 4.59e-21
C883 a_3368_n3928# a_3434_n4026# 3.89e-19
C884 a_3946_174# a_5360_46# 0.031298f
C885 a_5402_n1066# a_5456_n1194# 0.044963f
C886 B15 a_5773_n1814# 3.52e-21
C887 a_3589_n3928# a_3543_n2822# 0.001075f
C888 a_798_n1194# a_2273_n254# 2.74e-19
C889 a_894_n828# a_143_n1036# 2.9e-19
C890 a_n71_n4320# B4 8.21e-21
C891 a_4000_n3674# a_2995_n4294# 0.001187f
C892 a_3946_n1066# a_3946_n2306# 0.0016f
C893 a_3874_n1220# a_2995_n4294# 0.010503f
C894 a_3861_n600# a_4523_n574# 0.005159f
C895 a_3765_n600# a_4691_n574# 0.074717f
C896 a_3543_n342# a_6023_n574# 4.81e-19
C897 a_798_n3674# a_n131_n4294# 0.001991f
C898 a_3322_n4062# a_4000_n3308# 0.003825f
C899 a_4204_n3054# a_3904_n3674# 2.01e-19
C900 a_143_n2276# a_798_n3674# 1.17e-20
C901 B5 a_1201_n1814# 2.37e-19
C902 B6 B4 0.013937f
C903 B6 a_636_n3054# 9.78e-20
C904 a_2995_n4294# a_3946_174# 2.18e-19
C905 DVDD a_3627_n254# 2.46e-19
C906 a_636_n4294# a_1201_n3054# 1.04e-19
C907 a_101_n3674# a_1201_n4294# 0.003559f
C908 a_3736_n2068# a_4000_n2068# 1.31e-19
C909 a_3874_n1220# a_4204_n574# 0.026336f
C910 a_3543_n342# a_4523_n1814# 0.002766f
C911 a_3832_n2068# a_3904_n2434# 0.004869f
C912 a_3669_n342# a_3685_n1775# 2.79e-19
C913 a_3946_n1066# a_3322_n1582# 0.142863f
C914 A7 a_1997_n2434# 6.84e-21
C915 B14 a_5819_46# 8.1e-22
C916 B4 a_143_n3516# 0.002602f
C917 a_5773_n574# a_5855_n574# 0.006406f
C918 a_636_n3054# a_143_n3516# 0.102258f
C919 A11 a_3543_n2822# 0.004919f
C920 A13 a_3543_n342# 1.84e-20
C921 B1 a_2908_n600# 7.51e-21
C922 a_3946_174# a_4204_n574# 0.057421f
C923 a_143_n2276# a_1557_n1194# 0.018458f
C924 A9 a_4697_n2434# 5.03e-19
C925 a_2995_n4294# a_4523_n574# 1.89e-19
C926 a_2315_n4255# a_3322_n4062# 2.02e-20
C927 A10 B8 1.68e-19
C928 a_185_n3674# a_n131_n4294# 0.001149f
C929 a_1291_n1814# a_143_n1036# 1.59e-20
C930 DVDD a_1641_412# 0.160791f
C931 A6 a_n71_n4320# 0.081598f
C932 a_3832_n2434# a_4000_n2434# 2.18e-19
C933 A13 a_4441_n574# 0.076981f
C934 A7 a_2422_n3674# 7.66e-19
C935 a_n131_n3054# a_2315_n1775# 6e-20
C936 a_1201_n3054# a_1261_n1840# 5.51e-20
C937 A6 B6 1.27934f
C938 a_1557_n2434# a_2995_n4294# 0.004915f
C939 a_3322_n1582# a_4691_n574# 5.44e-19
C940 a_5819_n3674# a_4204_n3054# 0.033252f
C941 a_101_n2434# a_11_n2068# 0.006823f
C942 a_4204_n574# a_4523_n574# 0.003613f
C943 a_798_n2434# a_966_n2434# 0.00792f
C944 a_2908_n600# a_1641_n828# 5.23e-20
C945 B1 a_3874_20# 2.79e-20
C946 A1 a_3946_174# 2.18e-20
C947 a_636_n1814# a_894_n1194# 2.34e-19
C948 a_101_n1194# a_966_n1194# 3.46e-19
C949 DVDD a_n131_n1814# 1.03216f
C950 a_n71_n600# a_n131_n1814# 0.001041f
C951 a_143_n2276# a_1647_n574# 2.87e-19
C952 A6 a_143_n3516# 0.467991f
C953 Cin a_636_n574# 0.175088f
C954 A1 a_101_46# 1.36e-19
C955 a_3322_n1582# a_3368_n1775# 0.006879f
C956 A15 a_3861_n600# 3.72e-19
C957 A6 a_894_n3674# 5.43e-19
C958 a_5402_174# a_3543_n342# 2.69e-19
C959 B15 a_5360_n1194# 2.55e-19
C960 a_3434_n4026# B10 1.57e-20
C961 a_2273_n254# a_1201_n1814# 0.471487f
C962 a_3874_n1220# a_5402_n1066# 0.201352f
C963 B4 a_n131_n4294# 4.07e-19
C964 A3 a_2254_n1194# 0.114346f
C965 a_5819_n3308# a_5402_n3546# 0.030161f
C966 a_636_n1814# a_143_n1036# 0.026336f
C967 a_143_n2276# B4 0.674621f
C968 a_636_n3054# a_n131_n4294# 5.56e-19
C969 a_1557_n2434# a_1201_n4294# 0.016609f
C970 a_101_n1194# a_2273_n254# 5.68e-21
C971 a_3669_n2822# B10 4.1e-19
C972 a_143_n2276# a_636_n3054# 0.195149f
C973 a_3434_n1546# a_3669_n2822# 3.6e-19
C974 DVDD a_11_n3674# 2.33e-19
C975 B3 a_143_n1036# 0.020606f
C976 B0 a_185_n828# 5.74e-19
C977 Cin a_2422_n1194# 2.14e-20
C978 A0 a_541_n828# 3.08e-21
C979 DVDD a_798_n1194# 0.236555f
C980 B9 a_3946_n3546# 3.5e-19
C981 a_5402_174# a_4441_n574# 0.005909f
C982 a_5456_n3308# a_5819_n3308# 0.009846f
C983 a_1557_n1194# a_1968_n1814# 0.116264f
C984 A15 a_2995_n4294# 0.010491f
C985 a_3832_n1194# a_2908_n600# 0.005587f
C986 a_636_n3054# a_1641_n3308# 1.77e-21
C987 Cin a_2350_46# 4.74e-19
C988 A1 a_1997_46# 0.046632f
C989 DVDD a_2497_n4255# 8.63e-19
C990 a_315_n574# a_n131_n574# 0.00528f
C991 a_2995_n4294# B8 0.677478f
C992 a_143_n1036# a_1291_n574# 0.016475f
C993 a_5402_n2306# a_5288_n2068# 4.35e-21
C994 B2 a_894_n828# 2.91e-19
C995 A2 a_966_n828# 1.05e-19
C996 a_3832_n2434# a_3904_n2434# 0.005587f
C997 A10 a_5288_n3674# 5.43e-19
C998 A15 a_4204_n574# 0.011053f
C999 A6 a_n131_n4294# 0.02685f
C1000 S15 a_636_n574# 4.41e-21
C1001 A2 a_101_46# 0.003407f
C1002 A2 a_n71_n1840# 0.081598f
C1003 a_4204_n574# a_5819_n828# 0.091015f
C1004 a_541_n2434# a_n131_n1814# 0.001136f
C1005 a_1641_n2068# B5 0.020016f
C1006 A9 a_3434_n1546# 5.1e-20
C1007 DVDD a_315_n1814# 0.009564f
C1008 A11 a_3946_n3546# 0.791917f
C1009 a_2254_n2434# a_3874_n2460# 2.15e-20
C1010 a_1997_n3308# a_2995_n4294# 9.47e-19
C1011 a_3832_n2068# B9 2.91e-19
C1012 B1 a_636_n1814# 1.11e-19
C1013 a_1479_n1494# A3 0.001028f
C1014 A9 a_4363_n2434# 0.051667f
C1015 A7 a_1479_n3974# 0.001028f
C1016 a_3946_n2306# A5 2.18e-20
C1017 DVDD a_1997_n2434# 8.16e-19
C1018 a_3669_n2822# a_3711_n2734# 0.001239f
C1019 a_3765_n3080# a_3627_n2734# 3.31e-19
C1020 a_3434_n4026# a_5773_n4294# 1.26e-20
C1021 B2 a_n71_n3080# 2.27e-21
C1022 Cin B15 1.52e-20
C1023 DVDD A4 0.494087f
C1024 B1 B3 0.005115f
C1025 a_2783_n1775# a_2569_n1775# 0.005572f
C1026 A11 a_5360_n3674# 0.001236f
C1027 a_1557_n2434# a_2315_n1775# 9.88e-20
C1028 a_5773_n4294# a_3669_n2822# 3.93e-19
C1029 a_4441_n4294# a_3765_n3080# 7.34e-21
C1030 a_3655_n3996# a_3861_n3080# 5.6e-20
C1031 a_636_n3054# a_1968_n1814# 1.74e-20
C1032 a_4691_n1814# A9 7.81e-20
C1033 a_4691_n3054# a_3874_n3700# 1.21e-19
C1034 a_3543_n2822# a_5773_n3054# 0.001041f
C1035 a_3669_n2822# a_4441_n3054# 3.76e-19
C1036 a_3765_n3080# a_3861_n3080# 0.197466f
C1037 A14 a_5773_n3054# 1.82e-21
C1038 DVDD a_4691_n3054# 0.238543f
C1039 a_5192_n3674# a_5456_n3674# 8.12e-20
C1040 a_2254_n2434# a_n131_n3054# 3.5e-19
C1041 a_636_n574# a_966_46# 3.15e-19
C1042 a_1201_n574# a_2254_n1194# 4.56e-19
C1043 a_1201_n1814# a_1997_n828# 4.28e-19
C1044 B15 a_3669_n342# 0.081283f
C1045 a_2254_n3674# a_1201_n3054# 4.56e-19
C1046 a_1997_n3308# a_1201_n4294# 4.28e-19
C1047 a_1557_n1194# a_1467_n828# 0.006823f
C1048 DVDD a_185_n3308# 0.165024f
C1049 a_636_n1814# a_1641_n828# 0.12395f
C1050 B13 a_3832_46# 7.33e-20
C1051 A13 a_4000_46# 0.046632f
C1052 a_3655_n3996# a_3904_n2434# 7.07e-21
C1053 DVDD a_1201_n1814# 0.366096f
C1054 B3 a_1641_n828# 0.020016f
C1055 a_3765_n3080# a_3904_n2434# 4.74e-19
C1056 A5 a_1201_n3054# 0.081374f
C1057 a_101_n1194# a_n71_n600# 5.92e-19
C1058 DVDD a_101_n1194# 0.395339f
C1059 B1 a_1291_n574# 0.05645f
C1060 B10 a_6023_n4294# 0.056624f
C1061 a_315_n3054# a_n71_n3080# 0.006406f
C1062 a_1997_412# a_2350_412# 2.18e-19
C1063 a_5402_n1066# A15 1.36e-19
C1064 a_5288_412# a_5456_412# 2.18e-19
C1065 a_5402_n1066# a_5819_n828# 0.030161f
C1066 a_5402_n3546# B10 0.181244f
C1067 a_5402_n1066# B8 3.81e-20
C1068 a_2497_n4255# a_2569_n4255# 6.64e-19
C1069 B15 a_3874_n2460# 1.13e-19
C1070 a_2995_n4294# a_3861_n600# 0.001235f
C1071 A9 a_4441_n3054# 0.076981f
C1072 a_2995_n4294# a_1479_n2734# 1.25e-19
C1073 B2 a_636_n1814# 0.013754f
C1074 a_2254_n3674# a_636_n4294# 0.06247f
C1075 DVDD a_4441_n1814# 0.191496f
C1076 a_798_n2434# a_894_n2068# 0.004869f
C1077 a_541_n2068# a_966_n2068# 1.31e-19
C1078 a_1261_n4320# a_n131_n3054# 9.27e-21
C1079 a_5456_n3308# B10 0.017703f
C1080 B12 A14 1.68e-19
C1081 A12 B14 1.48e-19
C1082 a_101_46# a_636_n574# 0.172114f
C1083 B2 B3 0.003904f
C1084 a_3832_n828# a_3669_n342# 1.5e-20
C1085 a_4363_n828# a_2908_n600# 1.55e-19
C1086 A5 a_636_n4294# 0.004204f
C1087 a_5402_174# a_4000_46# 5.42e-21
C1088 Cin a_3177_n1814# 0.001873f
C1089 B11 a_4523_n4294# 0.007771f
C1090 a_541_n2434# A4 0.047225f
C1091 a_4691_n254# a_3765_n600# 0.004527f
C1092 A9 a_4000_n2068# 0.011819f
C1093 a_4204_n574# a_3861_n600# 0.182595f
C1094 a_4204_n574# a_5360_46# 0.0021f
C1095 a_4000_n3674# a_3904_n3674# 0.023012f
C1096 B13 a_4697_46# 6.45e-19
C1097 DVDD a_6023_n1814# 0.263219f
C1098 B11 a_1557_n3674# 2.32e-20
C1099 a_143_n3516# a_1201_n3054# 0.068052f
C1100 a_2273_n2734# a_n131_n3054# 0.158736f
C1101 a_2497_n1775# a_n131_n1814# 9.8e-19
C1102 a_147_n2734# a_n131_n4294# 6.93e-20
C1103 a_3946_n2306# a_5402_n2306# 0.003292f
C1104 a_6023_n254# a_5773_n574# 0.007234f
C1105 a_3874_20# a_4363_n828# 1.77e-21
C1106 B9 a_3832_n2434# 7.33e-20
C1107 a_636_n1814# a_1641_46# 1.55e-21
C1108 a_541_n2434# a_101_n1194# 4.36e-20
C1109 a_3322_n4062# a_4691_n4294# 1.57e-19
C1110 B6 a_966_n3308# 3.18e-19
C1111 a_1557_46# a_2459_n254# 3.34e-19
C1112 a_n71_n4320# a_636_n4294# 0.062036f
C1113 a_1261_n4320# a_101_n3674# 0.005934f
C1114 A5 a_1261_n1840# 9.85e-20
C1115 a_5773_n4294# a_6023_n4294# 0.025037f
C1116 B3 a_1641_46# 3.27e-20
C1117 a_2995_n4294# a_4204_n574# 0.00314f
C1118 a_5288_n3308# B10 2.91e-19
C1119 B14 a_3861_n3080# 2.57e-21
C1120 a_636_n574# a_1997_46# 0.045338f
C1121 B2 a_101_n2434# 5.99e-19
C1122 a_143_n3516# a_966_n3308# 2.69e-19
C1123 a_2273_n2734# a_894_n3308# 1.6e-20
C1124 B6 a_636_n4294# 0.013754f
C1125 a_3874_n3700# a_3322_n4062# 0.022847f
C1126 DVDD a_11_46# 2.33e-19
C1127 a_2569_n1448# a_3434_n1546# 3.16e-20
C1128 a_2995_n4294# a_1201_n4294# 0.008819f
C1129 a_3322_n1582# a_3736_n828# 1.91e-19
C1130 a_143_n2276# a_3946_n2306# 1.42e-20
C1131 B13 a_4441_n1814# 3.66e-21
C1132 a_5773_n4294# a_5402_n3546# 0.003994f
C1133 a_1467_n3674# a_798_n3674# 5.49e-20
C1134 DVDD a_3322_n4062# 1.15055f
C1135 Cin a_143_n1036# 0.043588f
C1136 a_636_n4294# a_143_n3516# 0.026336f
C1137 a_1261_n600# a_n131_n574# 0.041433f
C1138 A0 a_n131_n574# 0.025968f
C1139 a_2254_n2434# a_1557_n2434# 0.055111f
C1140 a_2350_n2068# a_636_n3054# 1.35e-20
C1141 a_101_n3674# a_2273_n2734# 5.68e-21
C1142 B5 a_1261_n3080# 0.214186f
C1143 DVDD a_1479_n3974# 5.64e-19
C1144 a_5360_n2434# a_5456_n2434# 0.023012f
C1145 a_894_n3674# a_636_n4294# 2.34e-19
C1146 a_5402_174# a_5192_46# 3.46e-19
C1147 a_966_n3674# a_101_n3674# 3.46e-19
C1148 a_3874_n1220# B15 1.25417f
C1149 B11 a_3736_n3308# 3.18e-19
C1150 a_5402_n1066# a_3861_n600# 2.05e-19
C1151 B4 a_n41_n3054# 0.056561f
C1152 a_636_n3054# a_n41_n3054# 4.33e-19
C1153 a_143_n2276# a_3322_n1582# 0.002815f
C1154 a_2273_n254# a_3543_n342# 4.14e-19
C1155 a_541_n2068# a_n131_n1814# 0.003779f
C1156 A14 a_5192_n1194# 7.66e-19
C1157 DVDD a_5288_n828# 4.94e-19
C1158 a_2995_n4294# a_1467_n3308# 5.92e-21
C1159 Cin a_2569_n1775# 0.089244f
C1160 a_1997_n3674# a_2422_n3674# 8.12e-20
C1161 a_5402_n1066# a_5360_46# 9.75e-22
C1162 B11 a_4363_n3308# 0.020016f
C1163 A14 a_3874_20# 4.45e-19
C1164 a_1201_n3054# a_n131_n4294# 6.83e-19
C1165 B15 a_3946_174# 4.05e-20
C1166 a_143_n2276# a_1201_n3054# 0.011525f
C1167 DVDD a_4697_n2068# 4.94e-19
C1168 B9 a_3765_n3080# 0.097286f
C1169 a_5402_174# a_5456_n828# 4.9e-19
C1170 a_1641_n2068# DVDD 0.160791f
C1171 a_1997_46# a_2350_46# 2.18e-19
C1172 a_3736_n2068# a_3322_n4062# 4.54e-21
C1173 a_3832_n3308# a_3322_n4062# 2.27e-19
C1174 a_2783_n4255# a_3543_n2822# 3.93e-20
C1175 a_5402_n1066# a_2995_n4294# 7.45e-19
C1176 A7 a_1261_n3080# 1.75e-19
C1177 a_3904_46# a_3832_46# 0.005587f
C1178 a_315_n574# a_n131_n1814# 2.52e-19
C1179 a_3861_n600# a_5855_n574# 0.00528f
C1180 A12 a_6153_412# 5.12e-20
C1181 B12 a_5819_412# 0.033026f
C1182 a_966_n3308# a_n131_n4294# 3.51e-20
C1183 a_4204_n3054# a_4363_n3308# 0.00341f
C1184 a_3322_n4062# a_4697_n3308# 1.07e-20
C1185 a_1557_n1194# B5 2.43e-20
C1186 a_3874_n1220# a_3832_n828# 1.35e-20
C1187 A6 a_n41_n3054# 7.55e-19
C1188 A0 a_541_412# 0.011819f
C1189 DVDD a_798_46# 0.236488f
C1190 B0 a_185_412# 0.033026f
C1191 a_636_n4294# a_n131_n4294# 0.044377f
C1192 Cin B1 0.091476f
C1193 a_143_n2276# a_636_n4294# 0.00167f
C1194 a_3226_n1582# a_3434_n1546# 0.190276f
C1195 a_5402_n1066# a_4204_n574# 0.219575f
C1196 A11 a_3655_n3996# 0.002825f
C1197 a_1557_n2434# a_2273_n2734# 0.008526f
C1198 A7 a_798_n3674# 0.001236f
C1199 A11 a_3765_n3080# 1.85e-19
C1200 a_2497_n1775# a_1201_n1814# 2.79e-19
C1201 A13 a_3765_n600# 0.081374f
C1202 B8 a_6023_n2734# 0.002402f
C1203 DVDD a_185_n2434# 0.003141f
C1204 a_143_n2276# a_3946_n1066# 1.4e-19
C1205 a_2569_n4255# a_3322_n4062# 2.95e-19
C1206 a_3322_n1582# a_1968_n1814# 1.71e-19
C1207 a_636_n4294# a_1641_n3308# 0.12395f
C1208 a_1997_n1194# a_2422_n1194# 8.12e-20
C1209 a_1997_n3308# a_2350_n3308# 2.18e-19
C1210 a_4000_n2434# a_4363_n2434# 0.008475f
C1211 a_5855_n3054# a_3543_n2822# 2.52e-19
C1212 a_4523_n3054# a_3765_n3080# 0.001897f
C1213 a_4691_n3054# a_3669_n2822# 2.26e-19
C1214 a_1997_n2068# A5 0.011819f
C1215 a_5360_n2434# A8 0.114467f
C1216 a_1201_n4294# a_2315_n1775# 3.16e-19
C1217 a_2254_n3674# A5 2.18e-20
C1218 a_143_n2276# a_1261_n1840# 0.015687f
C1219 a_2995_n4294# a_3685_n1775# 2.57e-19
C1220 a_4204_n574# a_5855_n574# 8.43e-19
C1221 a_143_n1036# a_966_46# 1.96e-19
C1222 a_2908_n600# a_2254_n1194# 0.004747f
C1223 a_1641_n1194# a_1201_n1814# 9.33e-19
C1224 a_541_n2068# A4 0.011819f
C1225 B4 B5 0.003904f
C1226 a_1557_n1194# a_966_n1194# 3.2e-20
C1227 a_636_n3054# B5 1.25937f
C1228 a_101_n1194# a_1641_n1194# 1.11e-20
C1229 DVDD a_3543_n342# 1.02027f
C1230 A15 B15 1.25275f
C1231 a_3322_n1582# a_4523_n1814# 3.9e-20
C1232 B3 a_1467_n1194# 6.45e-19
C1233 a_5402_174# a_3765_n600# 0.003561f
C1234 B1 S15 8.13e-22
C1235 a_2995_n4294# a_3368_n4255# 3.88e-19
C1236 A14 A8 0.00475f
C1237 A8 a_3543_n2822# 3.84e-19
C1238 A13 a_3322_n1582# 4.12e-19
C1239 A3 a_2422_n828# 1.05e-19
C1240 a_3861_n3080# B10 7.86e-19
C1241 a_143_n2276# a_3368_n1775# 0.001639f
C1242 a_1557_n1194# a_2273_n254# 0.142863f
C1243 DVDD a_4441_n574# 0.173165f
C1244 a_541_n2068# a_101_n1194# 1.79e-19
C1245 A2 a_185_n1194# 0.050725f
C1246 A9 a_4691_n3054# 0.007493f
C1247 a_3655_n1516# a_3765_n3080# 2.07e-19
C1248 A14 a_5773_n1814# 0.081598f
C1249 a_3434_n1546# a_3861_n3080# 4.03e-21
C1250 a_3322_n4062# a_3736_n2434# 2.27e-20
C1251 a_966_n828# a_143_n1036# 2.69e-19
C1252 a_541_n2434# a_185_n2434# 0.008475f
C1253 a_1557_46# a_n131_n574# 0.060379f
C1254 a_101_46# a_143_n1036# 0.008359f
C1255 a_143_n1036# a_n71_n1840# 1.52e-19
C1256 a_3736_n2068# a_3543_n342# 4.28e-20
C1257 a_1997_n2068# a_143_n3516# 1.25e-20
C1258 a_3832_n1194# a_3669_n342# 6.23e-20
C1259 a_3434_n1546# a_3904_n2434# 4.57e-19
C1260 a_2254_n3674# a_143_n3516# 2.01e-19
C1261 DVDD a_5819_n2434# 0.001386f
C1262 a_1997_n3308# a_2273_n2734# 0.003825f
C1263 a_2459_n254# a_1201_n574# 0.009339f
C1264 a_2363_n254# a_1201_n1814# 1.46e-22
C1265 DVDD a_4691_n3974# 4.62e-19
C1266 A1 a_1467_46# 5.03e-19
C1267 Cin a_1641_46# 0.002621f
C1268 a_2273_n254# a_1647_n574# 3.8e-19
C1269 A5 a_143_n3516# 0.051784f
C1270 a_2569_n1448# a_n131_n1814# 0.001075f
C1271 a_1557_n3674# a_n131_n3054# 6.4e-19
C1272 a_5360_n2434# a_4204_n3054# 0.002098f
C1273 B11 a_3543_n2822# 0.00432f
C1274 A10 a_5819_n3674# 0.050725f
C1275 B13 a_3543_n342# 2.07e-21
C1276 a_1261_n1840# a_1968_n1814# 0.053796f
C1277 DVDD a_1261_n3080# 0.17389f
C1278 B9 a_4697_n2434# 6.45e-19
C1279 A9 a_4441_n1814# 9.85e-20
C1280 DVDD a_1997_412# 0.154852f
C1281 a_5192_46# a_5456_46# 8.12e-20
C1282 a_2254_n2434# a_2995_n4294# 0.005482f
C1283 B6 a_n71_n4320# 0.226175f
C1284 a_2350_n3308# a_2995_n4294# 4.78e-20
C1285 A13 a_3946_n1066# 2.88e-19
C1286 a_3434_n4026# a_3322_n4062# 0.14976f
C1287 B13 a_4441_n574# 0.214186f
C1288 a_143_n1036# a_1997_46# 7.87e-20
C1289 B7 a_2422_n3674# 6.11e-20
C1290 A6 A7 0.019542f
C1291 a_5360_n2434# a_5192_n2068# 0.007578f
C1292 a_3669_n2822# a_3322_n4062# 0.471487f
C1293 a_3543_n2822# a_4204_n3054# 0.012648f
C1294 a_101_n2434# a_185_n2068# 0.030161f
C1295 a_3765_n3080# a_3795_n2734# 0.006083f
C1296 a_2995_n4294# a_3904_n3674# 0.009179f
C1297 a_5192_412# a_5360_46# 0.007578f
C1298 a_n71_n4320# a_143_n3516# 1.52e-19
C1299 a_3946_n2306# a_4000_n3308# 5.56e-19
C1300 a_3874_n2460# a_4363_n3308# 1.77e-21
C1301 B2 a_n131_n3054# 2.57e-21
C1302 DVDD a_798_n3674# 0.236555f
C1303 a_5773_n4294# a_3861_n3080# 1.01e-20
C1304 a_4441_n4294# a_4441_n3054# 0.002078f
C1305 a_101_n3674# a_1557_n3674# 0.003292f
C1306 B1 a_3946_174# 2.32e-20
C1307 a_3736_n1194# a_3322_n1582# 4.57e-19
C1308 B6 a_143_n3516# 0.662565f
C1309 A0 a_n131_n1814# 3.84e-19
C1310 a_3765_n3080# a_5773_n3054# 2.84e-19
C1311 a_3861_n3080# a_4441_n3054# 0.041433f
C1312 A1 a_636_n574# 0.512147f
C1313 B1 a_101_46# 7.19e-19
C1314 DVDD a_6023_n3054# 0.242051f
C1315 a_2254_n2434# a_1201_n4294# 3.97e-19
C1316 a_1201_n1814# a_2350_n828# 1.5e-20
C1317 B6 a_894_n3674# 7.33e-20
C1318 a_2350_n3308# a_1201_n4294# 1.5e-20
C1319 a_2254_n3674# a_n131_n4294# 0.008425f
C1320 B15 a_3861_n600# 8.88e-19
C1321 a_1997_n2068# a_143_n2276# 0.012702f
C1322 a_1557_n1194# a_1997_n828# 0.004914f
C1323 a_636_n1814# a_2254_n1194# 0.06247f
C1324 a_2254_n3674# a_143_n2276# 0.003114f
C1325 a_2350_n1194# a_143_n2276# 1.22e-19
C1326 A14 a_5360_n1194# 0.114467f
C1327 A5 a_n131_n4294# 1.84e-20
C1328 A13 a_4691_n574# 0.007493f
C1329 B3 a_2254_n1194# 0.077341f
C1330 a_143_n2276# A5 0.060612f
C1331 DVDD a_1557_n1194# 0.387599f
C1332 a_315_n3054# a_n131_n3054# 0.00528f
C1333 a_1291_n3054# a_1261_n3080# 0.025037f
C1334 a_894_n3674# a_143_n3516# 1.28e-19
C1335 a_1261_n4320# a_2995_n4294# 8.92e-19
C1336 DVDD a_185_n3674# 0.003788f
C1337 A0 a_798_n1194# 2.18e-20
C1338 Cin a_185_n828# 1.77e-21
C1339 A3 a_n131_n574# 3.72e-19
C1340 a_541_n3674# a_966_n3674# 8.12e-20
C1341 a_3226_n1582# a_n131_n1814# 7.26e-19
C1342 A9 a_3322_n4062# 4.12e-19
C1343 a_4204_n574# a_5192_412# 2.91e-20
C1344 A13 a_2254_46# 9.68e-20
C1345 a_3904_n2434# a_4000_n2068# 0.02283f
C1346 a_5456_n3674# a_5402_n2306# 4.36e-20
C1347 DVDD a_6153_n1194# 2.33e-19
C1348 B15 a_2995_n4294# 0.010735f
C1349 A5 a_1641_n3308# 1.58e-21
C1350 a_2995_n4294# a_2273_n2734# 0.025133f
C1351 A1 a_2350_46# 5.43e-19
C1352 Cin a_2422_46# 5.78e-19
C1353 DVDD a_4000_46# 8.16e-19
C1354 B1 a_1997_46# 0.005557f
C1355 a_5360_n3674# A8 2.18e-20
C1356 DVDD a_147_n1494# 0.001263f
C1357 a_1261_n4320# a_1201_n4294# 0.188936f
C1358 a_n71_n4320# a_n131_n4294# 0.188784f
C1359 a_1968_n4294# a_n131_n3054# 5.85e-21
C1360 a_5855_n1814# B14 0.007771f
C1361 a_2315_n4255# a_1201_n3054# 2.4e-19
C1362 a_4363_n828# a_3669_n342# 3.93e-19
C1363 a_5192_n828# a_2908_n600# 4.71e-21
C1364 B2 a_966_n828# 3.18e-19
C1365 DVDD a_1647_n574# 0.005567f
C1366 B15 a_4204_n574# 0.020606f
C1367 A2 a_11_n1194# 4.78e-19
C1368 a_966_n2434# A4 7.66e-19
C1369 a_1997_n1194# a_143_n1036# 4.76e-20
C1370 B6 a_n131_n4294# 0.057188f
C1371 B2 a_101_46# 1.3e-19
C1372 a_6023_n254# a_3861_n600# 0.002789f
C1373 A2 a_636_n574# 4.45e-19
C1374 a_1557_n2434# a_1557_n3674# 0.007318f
C1375 B2 a_n71_n1840# 0.226175f
C1376 a_3322_n1582# a_3832_412# 1.21e-20
C1377 B9 a_3434_n1546# 0.001196f
C1378 DVDD a_4691_n1494# 4.62e-19
C1379 a_2569_n1448# a_1201_n1814# 6.39e-19
C1380 DVDD B4 0.801352f
C1381 DVDD a_636_n3054# 0.915951f
C1382 B11 a_3946_n3546# 0.175017f
C1383 a_2273_n2734# a_1201_n4294# 0.471487f
C1384 a_2363_n2734# a_1201_n3054# 0.006083f
C1385 a_3589_n1448# a_3669_n342# 6.39e-19
C1386 a_5456_n2068# a_3543_n342# 0.003779f
C1387 a_143_n3516# a_n131_n4294# 0.012648f
C1388 a_143_n2276# a_143_n3516# 0.045171f
C1389 a_2254_n2434# a_2315_n1775# 4e-19
C1390 a_894_n3674# a_n131_n4294# 1.41e-19
C1391 a_2254_n3674# a_1968_n1814# 4.29e-21
C1392 a_1479_n1494# B3 0.002951f
C1393 B9 a_4363_n2434# 0.019568f
C1394 B7 a_1479_n3974# 0.002951f
C1395 a_3946_n2306# B5 2.32e-20
C1396 a_2995_n4294# a_3832_n828# 2.35e-20
C1397 A2 a_11_n828# 5.12e-20
C1398 a_1968_n4294# a_101_n3674# 4.58e-20
C1399 a_2315_n4255# a_636_n4294# 9.72e-19
C1400 A5 a_1968_n1814# 5.1e-20
C1401 B11 a_5360_n3674# 2.55e-19
C1402 a_4691_n1814# B9 2.83e-19
C1403 B14 a_5773_n3054# 2.27e-21
C1404 a_2273_n2734# a_1467_n3308# 1.07e-20
C1405 a_5402_n3546# a_3322_n4062# 5.68e-21
C1406 a_3946_n3546# a_4204_n3054# 0.005791f
C1407 a_143_n3516# a_1641_n3308# 0.00341f
C1408 a_101_46# a_1641_46# 1.11e-20
C1409 a_3322_n1582# a_4000_n828# 0.003825f
C1410 A14 a_3669_n342# 1.6e-19
C1411 a_3669_n2822# a_3543_n342# 1.08e-20
C1412 a_4204_n574# a_3832_n828# 1.19e-20
C1413 A11 B10 1.74e-19
C1414 B13 a_4000_46# 0.005557f
C1415 a_3177_n1814# a_2995_n4294# 0.00462f
C1416 a_5360_n2434# a_3874_n2460# 0.012687f
C1417 B5 a_1201_n3054# 0.097286f
C1418 a_n131_n574# a_1201_n574# 0.197466f
C1419 a_1261_n600# a_1201_n1814# 3.76e-19
C1420 DVDD A6 0.502539f
C1421 a_1557_46# a_1641_412# 0.030161f
C1422 A0 a_101_n1194# 6.66e-20
C1423 a_5360_n3674# a_4204_n3054# 0.079554f
C1424 a_1641_n3674# a_101_n3674# 1.11e-20
C1425 a_1997_412# a_2422_412# 1.31e-19
C1426 a_2254_46# a_2350_412# 0.004869f
C1427 a_5402_n1066# B15 7.19e-19
C1428 A14 a_5773_n574# 0.001913f
C1429 a_5360_46# a_5456_412# 0.02283f
C1430 a_2273_n254# a_3765_n600# 2.76e-20
C1431 A11 a_4363_n2434# 1.4e-21
C1432 a_636_n3054# a_1291_n3054# 0.006212f
C1433 A14 a_5456_n1194# 0.047225f
C1434 a_894_n2068# a_n131_n1814# 2.73e-20
C1435 DVDD a_5456_n828# 0.1561f
C1436 DVDD a_5288_n2068# 4.94e-19
C1437 a_3874_n2460# a_3543_n2822# 5.56e-19
C1438 a_143_n2276# a_n131_n4294# 0.525748f
C1439 a_541_n2434# B4 0.005557f
C1440 a_894_n2434# a_101_n2434# 3.78e-19
C1441 B9 a_4441_n3054# 0.214186f
C1442 a_1557_46# a_n131_n1814# 7.63e-19
C1443 a_4691_n3974# a_3434_n4026# 3.05e-19
C1444 a_1641_46# a_1997_46# 0.008475f
C1445 A9 a_3543_n342# 8.47e-19
C1446 a_2273_n2734# a_2315_n1775# 8.08e-22
C1447 B12 B14 0.013937f
C1448 a_1997_n3308# a_1557_n3674# 0.004914f
C1449 a_2569_n3928# a_2995_n4294# 3.4e-19
C1450 a_4691_n3974# a_3669_n2822# 0.002666f
C1451 B5 a_636_n4294# 1.11e-19
C1452 a_6023_n3974# a_3543_n2822# 0.002687f
C1453 a_2543_n254# a_n131_n1814# 2.77e-20
C1454 A7 a_1201_n3054# 1.85e-19
C1455 B9 a_4000_n2068# 0.005326f
C1456 a_1968_n4294# a_1557_n2434# 2.72e-21
C1457 a_3322_n4062# a_5288_n3308# 1.6e-20
C1458 a_4204_n3054# a_5192_n3308# 2.69e-19
C1459 a_143_n2276# a_1641_n3308# 4.14e-19
C1460 a_541_n828# a_894_n828# 2.18e-19
C1461 a_3832_n1194# A15 5.43e-19
C1462 a_3543_n2822# a_n131_n3054# 8.62e-20
C1463 a_3946_n1066# a_4000_n828# 0.004914f
C1464 a_3874_n1220# a_4363_n828# 0.12395f
C1465 a_143_n2276# a_541_n1194# 7.7e-21
C1466 a_3434_n1546# a_3655_n1516# 0.153192f
C1467 a_3322_n1582# a_2273_n254# 0.00968f
C1468 A11 a_5773_n4294# 1.38e-21
C1469 a_2569_n3928# a_1201_n4294# 6.39e-19
C1470 a_1557_n2434# a_2459_n2734# 3.34e-19
C1471 A6 a_541_n2434# 2.43e-21
C1472 A11 a_4441_n3054# 1.75e-19
C1473 B5 a_1261_n1840# 7.54e-19
C1474 a_2273_n254# a_1201_n3054# 4.56e-21
C1475 a_143_n2276# a_1479_n254# 1.26e-19
C1476 A7 a_636_n4294# 0.51166f
C1477 a_1997_n2068# a_2350_n2068# 2.18e-19
C1478 A0 a_11_46# 4.78e-19
C1479 Cin a_2254_n1194# 0.002539f
C1480 a_4441_n4294# a_4691_n3054# 9.75e-20
C1481 B14 a_2908_n600# 2.15e-21
C1482 a_2254_n3674# a_2422_n3308# 0.007578f
C1483 a_4523_n3054# a_4441_n3054# 0.006406f
C1484 a_4691_n3054# a_3861_n3080# 0.058037f
C1485 a_5819_n2068# A8 0.011602f
C1486 B0 a_n131_n574# 0.059236f
C1487 A1 a_143_n1036# 0.051784f
C1488 a_n131_n4294# a_1968_n1814# 1.28e-20
C1489 a_143_n2276# a_1968_n1814# 0.025299f
C1490 a_5192_n3674# a_3874_n3700# 3.15e-19
C1491 a_2908_n600# a_2422_n828# 2.11e-20
C1492 a_4697_n3674# a_3946_n3546# 0.006958f
C1493 a_101_n1194# a_541_46# 1.67e-20
C1494 a_5402_174# a_5288_46# 3.78e-19
C1495 a_5402_n3546# a_3543_n342# 2.04e-19
C1496 a_1557_n2434# a_2422_n2434# 3.12e-19
C1497 a_3832_n3674# a_3669_n2822# 6.23e-20
C1498 a_3874_n1220# A14 0.020957f
C1499 a_1557_n1194# a_1641_n1194# 0.06777f
C1500 a_185_n1194# a_143_n1036# 0.033252f
C1501 DVDD a_3765_n600# 0.179937f
C1502 DVDD a_147_n2734# 6.9e-19
C1503 B14 a_5192_n1194# 6.11e-20
C1504 B14 a_3874_20# 9.78e-20
C1505 a_5360_n3674# a_4697_n3674# 5.49e-20
C1506 a_5456_n3308# a_3543_n342# 2.21e-19
C1507 a_2995_n4294# a_4523_n4294# 1.4e-19
C1508 A3 a_n131_n1814# 0.004919f
C1509 A13 a_4691_n254# 9.63e-19
C1510 A8 a_3765_n3080# 4.94e-20
C1511 a_1997_46# a_2422_46# 8.12e-20
C1512 a_3946_n1066# a_2273_n254# 8.35e-21
C1513 a_143_n2276# a_4523_n1814# 1.35e-19
C1514 a_5773_n3054# B10 0.001373f
C1515 a_2254_n3674# a_2315_n4255# 6.53e-19
C1516 a_147_n254# a_n71_n600# 0.007234f
C1517 DVDD a_147_n254# 6.9e-19
C1518 A2 a_894_n1194# 5.43e-19
C1519 DVDD a_5819_n1194# 0.001386f
C1520 a_2995_n4294# a_1557_n3674# 0.005131f
C1521 a_3946_n2306# a_3874_n3700# 0.002601f
C1522 a_3874_20# a_4363_46# 0.033252f
C1523 a_n71_n4320# a_n41_n3054# 3.47e-20
C1524 B7 a_1261_n3080# 7.54e-19
C1525 a_1557_46# a_1201_n1814# 0.016609f
C1526 DVDD a_3946_n2306# 0.369711f
C1527 a_3904_46# a_4000_46# 0.023012f
C1528 a_798_n1194# A3 0.001236f
C1529 a_2273_n254# a_1261_n1840# 6.23e-19
C1530 a_2254_n2434# a_2273_n2734# 2.77e-19
C1531 B6 a_n41_n3054# 3.35e-19
C1532 a_2543_n254# a_1201_n1814# 0.008516f
C1533 a_2350_n3308# a_2273_n2734# 2.27e-19
C1534 a_3627_n254# a_1201_n574# 1.71e-20
C1535 A2 a_143_n1036# 0.467991f
C1536 DVDD a_894_412# 5.34e-19
C1537 B0 a_541_412# 0.017703f
C1538 A0 a_798_46# 0.114467f
C1539 Cin a_185_412# 0.090852f
C1540 A1 B1 1.25311f
C1541 A14 a_6023_n1494# 0.001052f
C1542 A15 a_4363_n828# 0.011964f
C1543 a_636_n3054# a_1641_n1194# 1.55e-21
C1544 a_n131_n3054# a_2254_n1194# 4.82e-21
C1545 DVDD a_3322_n1582# 1.15917f
C1546 B11 a_3655_n3996# 2.1e-19
C1547 a_n41_n1814# a_n131_n1814# 0.096176f
C1548 a_1557_n3674# a_1201_n4294# 0.044539f
C1549 a_143_n3516# a_n41_n3054# 0.002038f
C1550 a_143_n2276# a_1467_n828# 1.22e-20
C1551 B7 a_798_n3674# 2.55e-19
C1552 a_5360_n1194# a_5192_n828# 0.007578f
C1553 B11 a_3765_n3080# 0.00216f
C1554 B13 a_3765_n600# 0.097286f
C1555 DVDD a_1201_n3054# 0.180057f
C1556 a_2273_n254# a_2254_46# 2.77e-19
C1557 A1 a_1641_n828# 1.58e-21
C1558 a_2422_n2068# a_2995_n4294# 4.91e-20
C1559 a_3832_n2068# a_3874_n2460# 1.35e-20
C1560 a_541_n2068# B4 0.017703f
C1561 a_3627_n2734# a_3322_n4062# 7.04e-19
C1562 a_798_n2434# a_101_n2434# 0.057766f
C1563 a_3832_n1194# a_2995_n4294# 7.92e-20
C1564 a_3736_n3308# a_2995_n4294# 1.14e-19
C1565 a_4441_n4294# a_3322_n4062# 6.23e-19
C1566 a_5360_n2434# B8 0.078639f
C1567 a_1997_n2068# B5 0.005326f
C1568 a_1557_n3674# a_1467_n3308# 0.006823f
C1569 a_5456_n2068# a_5288_n2068# 2.18e-19
C1570 a_143_n1036# a_1467_46# 9.38e-21
C1571 a_1261_n4320# a_2273_n2734# 6.23e-19
C1572 a_3765_n3080# a_4204_n3054# 0.068052f
C1573 a_3861_n3080# a_3322_n4062# 0.158736f
C1574 a_2995_n4294# a_4363_n3308# 0.001123f
C1575 A5 a_2350_n2434# 5.43e-19
C1576 DVDD a_966_n3308# 7.01e-19
C1577 A5 B5 1.25311f
C1578 a_5773_n4294# a_5773_n3054# 0.001197f
C1579 a_4000_n1194# a_3322_n1582# 0.001323f
C1580 a_636_n3054# A9 2.02e-20
C1581 a_636_n4294# a_3874_n3700# 0.001289f
C1582 a_n131_n574# a_2908_n600# 3.32e-19
C1583 a_1201_n574# a_n131_n1814# 6.83e-19
C1584 DVDD a_636_n4294# 1.04604f
C1585 A15 A14 0.019542f
C1586 a_3322_n4062# a_3904_n2434# 2.77e-19
C1587 a_2350_n2068# a_143_n2276# 3.84e-19
C1588 a_2422_n3308# a_143_n2276# 4.05e-20
C1589 a_1557_n1194# a_2350_n828# 4.35e-21
C1590 a_3874_n1220# a_2254_n1194# 2.34e-21
C1591 a_4000_n3674# a_3946_n3546# 0.046215f
C1592 a_4363_n3674# a_3874_n3700# 0.033252f
C1593 A14 a_5819_n828# 0.011602f
C1594 B14 A8 1.23e-19
C1595 A14 B8 1.32e-19
C1596 B13 a_3322_n1582# 0.001085f
C1597 B8 a_3543_n2822# 4.07e-19
C1598 DVDD a_4363_n3674# 0.001386f
C1599 B3 a_2422_n828# 3.18e-19
C1600 DVDD a_3946_n1066# 0.387599f
C1601 a_1291_n3054# a_1201_n3054# 0.074717f
C1602 a_n41_n3054# a_n131_n4294# 4.81e-19
C1603 a_1647_n3054# a_n131_n3054# 0.005159f
C1604 a_1968_n4294# a_2995_n4294# 0.008558f
C1605 a_143_n2276# a_n41_n3054# 1.35e-19
C1606 B2 a_185_n1194# 0.021045f
C1607 B14 a_5773_n1814# 0.226175f
C1608 B9 a_4691_n3054# 0.05645f
C1609 A3 a_1201_n1814# 0.077871f
C1610 A10 a_5360_n2434# 1.29e-20
C1611 a_101_n1194# A3 1.36e-19
C1612 A7 a_2254_n3674# 0.114346f
C1613 a_5402_174# a_6153_46# 0.006958f
C1614 a_3434_n1546# a_2908_n600# 3.31e-19
C1615 a_3226_n1582# a_3543_n342# 0.015565f
C1616 a_4000_n2068# a_4363_n2068# 0.009846f
C1617 a_636_n574# a_143_n1036# 0.102258f
C1618 DVDD a_1261_n1840# 0.191496f
C1619 A7 A5 0.002462f
C1620 a_2995_n4294# a_2459_n2734# 2.17e-19
C1621 a_n41_n1814# A4 7.55e-19
C1622 a_5819_n3308# A8 7.78e-19
C1623 a_541_46# a_798_46# 0.023012f
C1624 a_2315_n4255# a_n131_n4294# 0.011237f
C1625 B15 a_3832_n828# 2.91e-19
C1626 a_1968_n4294# a_1201_n4294# 0.055436f
C1627 A1 a_1641_46# 0.051667f
C1628 B1 a_1467_46# 6.45e-19
C1629 a_1641_n3674# a_2995_n4294# 4.99e-19
C1630 B5 a_143_n3516# 0.046267f
C1631 a_143_n2276# a_2315_n4255# 0.040089f
C1632 DVDD a_4691_n574# 0.238543f
C1633 a_1641_n2434# a_1997_n2434# 0.008475f
C1634 a_636_n4294# a_1291_n3054# 1.21e-19
C1635 A10 a_3543_n2822# 0.02685f
C1636 A12 a_3543_n342# 3.84e-19
C1637 a_4000_n1194# a_3946_n1066# 0.046215f
C1638 a_11_n828# a_143_n1036# 1.23e-20
C1639 a_2350_n1194# a_2273_n254# 4.97e-19
C1640 a_2254_n3674# a_2273_n254# 5.66e-21
C1641 a_1557_n2434# a_2254_n1194# 9.75e-22
C1642 B9 a_4441_n1814# 7.54e-19
C1643 A11 a_4691_n3054# 7.81e-20
C1644 a_n41_n1814# a_1201_n1814# 2.66e-19
C1645 A2 B2 1.27934f
C1646 DVDD a_2254_46# 0.247054f
C1647 a_5288_46# a_5456_46# 2.18e-19
C1648 A5 a_2273_n254# 5.52e-19
C1649 DVDD a_3368_n1775# 0.001765f
C1650 A7 a_n71_n4320# 1.38e-21
C1651 a_2459_n2734# a_1201_n4294# 0.001239f
C1652 a_6153_n2068# a_3543_n342# 3.89e-20
C1653 a_143_n2276# a_2363_n2734# 0.00102f
C1654 B13 a_3946_n1066# 3.5e-19
C1655 A12 a_4441_n574# 6.77e-21
C1656 a_3946_n2306# a_3736_n2434# 3.12e-19
C1657 a_2995_n4294# a_2422_n2434# 1.79e-19
C1658 a_1641_n3674# a_1201_n4294# 9.33e-19
C1659 B6 A7 1.74e-19
C1660 A6 B7 2.69e-19
C1661 a_2995_n4294# a_4363_n828# 6.21e-19
C1662 a_5192_412# a_5456_412# 1.31e-19
C1663 a_1557_46# a_798_46# 0.031298f
C1664 A13 a_5402_174# 1.36e-19
C1665 a_3736_n828# a_4000_n828# 1.31e-19
C1666 A7 a_143_n3516# 0.011053f
C1667 a_101_46# a_185_412# 0.030161f
C1668 B0 a_n131_n1814# 4.07e-19
C1669 B1 a_636_n574# 1.25937f
C1670 a_5288_n3674# a_3543_n2822# 1.41e-19
C1671 A14 a_3861_n600# 2.3e-19
C1672 a_3861_n3080# a_3543_n342# 0.001229f
C1673 a_3765_n3080# a_3669_n342# 3.32e-21
C1674 a_3322_n1582# a_4697_n828# 1.07e-20
C1675 a_4204_n574# a_4363_n828# 0.00341f
C1676 a_3589_n1448# a_2995_n4294# 2.7e-19
C1677 a_5360_n2434# a_2995_n4294# 0.101686f
C1678 B14 a_5360_n1194# 0.078521f
C1679 a_143_n2276# a_2350_n2434# 6.26e-19
C1680 a_3904_46# a_3765_n600# 4.74e-19
C1681 B13 a_4691_n574# 0.05645f
C1682 A14 a_5360_46# 1.29e-20
C1683 a_1201_n574# a_1201_n1814# 0.15552f
C1684 A15 a_2254_n1194# 9.68e-20
C1685 B5 a_n131_n4294# 2.07e-21
C1686 a_143_n2276# B5 0.107685f
C1687 a_1557_n1194# a_1261_n600# 1.81e-19
C1688 a_636_n1814# a_n131_n574# 0.003854f
C1689 a_5819_n3308# a_4204_n3054# 0.091015f
C1690 a_1997_n3674# a_636_n4294# 0.045338f
C1691 a_3543_n342# a_3904_n2434# 0.002327f
C1692 a_636_n574# a_1641_n828# 1.77e-21
C1693 B0 a_798_n1194# 1.17e-20
C1694 Cin a_541_n828# 6.58e-21
C1695 B3 a_n131_n574# 8.88e-19
C1696 a_1467_n2068# a_n131_n1814# 3.89e-20
C1697 a_5360_n2434# a_4204_n574# 1.17e-20
C1698 B9 a_3322_n4062# 0.001085f
C1699 B13 a_2254_46# 1.77e-20
C1700 a_3434_n4026# a_3946_n2306# 2.72e-21
C1701 DVDD a_6153_n828# 5.28e-19
C1702 a_4204_n3054# a_4697_n2434# 9.38e-21
C1703 a_3946_n2306# a_3669_n2822# 0.016609f
C1704 A14 a_2995_n4294# 2.56e-19
C1705 a_3874_n2460# a_3765_n3080# 0.104793f
C1706 a_2995_n4294# a_3543_n2822# 0.542682f
C1707 a_966_n2434# B4 6.11e-20
C1708 a_966_n2434# a_636_n3054# 3.15e-19
C1709 Cin a_2459_n254# 5.54e-19
C1710 B5 a_1641_n3308# 9.06e-20
C1711 a_5360_n3674# B8 1.17e-20
C1712 B1 a_2350_46# 7.33e-20
C1713 A1 a_2422_46# 7.66e-19
C1714 a_4691_n3974# a_4441_n4294# 0.007234f
C1715 a_1997_n1194# a_2254_n1194# 0.023012f
C1716 a_2254_n2434# a_1557_n3674# 3.32e-21
C1717 a_n131_n574# a_1291_n574# 0.058037f
C1718 a_1261_n600# a_1647_n574# 0.006406f
C1719 a_2350_n3308# a_1557_n3674# 4.35e-21
C1720 a_2254_n3674# a_3874_n3700# 2.15e-20
C1721 a_1641_n2068# A3 1.58e-21
C1722 B2 a_11_n1194# 3.15e-19
C1723 a_3322_n1582# a_3669_n2822# 1.12e-20
C1724 A14 a_4204_n574# 0.467991f
C1725 DVDD a_1997_n2068# 0.154852f
C1726 B2 a_636_n574# 9.78e-20
C1727 A7 a_n131_n4294# 0.004919f
C1728 A7 a_143_n2276# 0.00207f
C1729 DVDD a_2254_n3674# 0.247054f
C1730 A8 B10 1.48e-19
C1731 a_1557_n3674# a_3904_n3674# 2.97e-20
C1732 a_3322_n1582# a_3904_46# 2.77e-19
C1733 a_3669_n2822# a_1201_n3054# 6.3e-20
C1734 a_3543_n2822# a_1201_n4294# 1.68e-20
C1735 a_3765_n3080# a_n131_n3054# 4.08e-20
C1736 DVDD A5 0.460573f
C1737 a_3946_n1066# a_4697_n828# 0.006823f
C1738 A10 a_3946_n3546# 0.001406f
C1739 A11 a_3322_n4062# 0.037805f
C1740 a_3434_n1546# a_5773_n1814# 1.26e-20
C1741 a_3946_n2306# A9 0.792469f
C1742 a_n41_n4294# a_1201_n4294# 2.66e-19
C1743 a_143_n2276# a_2790_n3928# 8.05e-19
C1744 A7 a_1641_n3308# 0.011964f
C1745 A2 a_185_n828# 0.011602f
C1746 B5 a_1968_n1814# 0.001196f
C1747 a_2273_n254# a_n131_n4294# 3.04e-20
C1748 A10 a_5360_n3674# 0.114467f
C1749 a_143_n2276# a_2273_n254# 0.039688f
C1750 a_5360_n2434# a_5402_n1066# 1.25e-21
C1751 a_4523_n3054# a_3322_n4062# 3.8e-19
C1752 a_1261_n4320# a_1557_n3674# 0.003171f
C1753 a_2254_n2434# a_2422_n2068# 0.007578f
C1754 a_636_n574# a_1641_46# 0.033252f
C1755 Cin a_2422_n828# 1.87e-20
C1756 B14 a_3669_n342# 4.1e-19
C1757 a_541_n1194# a_966_n1194# 8.12e-20
C1758 A9 a_3322_n1582# 5.52e-19
C1759 DVDD a_n71_n4320# 0.188115f
C1760 B11 B10 0.003904f
C1761 a_636_n4294# a_3669_n2822# 8.93e-21
C1762 a_6023_n3054# a_3861_n3080# 0.131556f
C1763 a_n131_n1814# a_2908_n600# 0.017585f
C1764 B0 a_101_n1194# 6.9e-19
C1765 DVDD B6 0.814551f
C1766 a_3368_n1448# a_1968_n1814# 8.12e-20
C1767 a_3177_n1814# a_2569_n1775# 7.45e-19
C1768 a_1557_46# a_1997_412# 0.004411f
C1769 a_3736_n3308# a_3904_n3674# 0.007578f
C1770 a_5192_n3674# a_5402_n3546# 3.46e-19
C1771 a_2254_46# a_2422_412# 0.007578f
C1772 a_1557_n3674# a_2273_n2734# 0.142863f
C1773 a_4363_n3674# a_3669_n2822# 9.33e-19
C1774 a_5402_n1066# A14 0.780011f
C1775 a_315_n4294# a_636_n4294# 8e-20
C1776 B14 a_5773_n574# 0.001373f
C1777 DVDD a_5456_n3674# 8.16e-19
C1778 a_894_n1194# a_143_n1036# 1.28e-19
C1779 A5 a_1291_n3054# 0.007493f
C1780 B11 a_4363_n2434# 3.27e-20
C1781 B14 a_5456_n1194# 0.005557f
C1782 DVDD a_143_n3516# 0.789008f
C1783 a_966_n3674# a_1557_n3674# 3.2e-20
C1784 a_3946_n1066# a_3904_46# 3.32e-21
C1785 a_798_n2434# a_101_n3674# 9.75e-22
C1786 A13 a_4000_n828# 8.69e-21
C1787 a_4204_n3054# B10 0.662565f
C1788 A10 a_5192_n3308# 1.05e-19
C1789 a_5360_n3674# a_5288_n3674# 0.005587f
C1790 a_5773_n4294# A8 2.8e-21
C1791 DVDD a_894_n3674# 8.89e-20
C1792 a_6153_n3308# a_3543_n342# 4.61e-21
C1793 a_894_n828# a_n131_n1814# 3.32e-20
C1794 A3 a_3543_n342# 9.21e-20
C1795 a_3655_n1516# a_3322_n4062# 8.08e-22
C1796 A8 a_4441_n3054# 6.77e-21
C1797 a_11_n2434# a_101_n2434# 0.006958f
C1798 B9 a_3543_n342# 7.3e-19
C1799 a_2995_n4294# a_3946_n3546# 0.007758f
C1800 a_4204_n3054# a_4363_n2434# 8.74e-19
C1801 B7 a_1201_n3054# 0.00216f
C1802 DVDD a_5402_n2306# 0.389244f
C1803 a_1557_n1194# a_1557_46# 0.007318f
C1804 a_1557_n2434# a_2543_n2734# 3.01e-19
C1805 a_3946_n1066# A9 1.91e-19
C1806 a_2273_n254# a_1968_n1814# 0.14976f
C1807 a_798_n1194# a_894_n828# 0.004869f
C1808 a_3832_n1194# B15 7.33e-20
C1809 a_541_n828# a_966_n828# 1.31e-19
C1810 Cin a_2790_n1448# 8.05e-19
C1811 a_2422_n2068# a_2273_n2734# 4.54e-21
C1812 A12 a_5192_46# 7.66e-19
C1813 a_5360_n3674# a_2995_n4294# 1.17e-20
C1814 DVDD a_3736_n828# 6.64e-19
C1815 a_n131_n1814# a_n71_n3080# 0.001891f
C1816 a_541_n828# a_101_46# 4.9e-19
C1817 a_6023_n1814# a_5773_n3054# 3.47e-20
C1818 a_2254_n3674# a_1997_n3674# 0.023012f
C1819 a_1291_n1814# a_n131_n1814# 0.017157f
C1820 B11 a_5773_n4294# 3.52e-21
C1821 a_143_n2276# a_1997_n828# 9.96e-19
C1822 a_143_n3516# a_1291_n3054# 0.016475f
C1823 a_3874_n3700# a_n131_n4294# 1.07e-20
C1824 a_3946_n3546# a_1201_n4294# 9.92e-21
C1825 a_3904_46# a_2254_46# 0.004465f
C1826 a_143_n2276# a_3874_n3700# 1.28e-20
C1827 A2 a_185_n2068# 6.72e-19
C1828 B11 a_4441_n3054# 7.54e-19
C1829 a_3946_174# a_3736_46# 3.12e-19
C1830 a_1261_n4320# a_1968_n4294# 0.053796f
C1831 DVDD a_n131_n4294# 0.916407f
C1832 A12 a_5456_n828# 3.08e-21
C1833 DVDD a_143_n2276# 1.81134f
C1834 a_636_n3054# a_3904_n2434# 2.15e-20
C1835 a_541_n2434# a_143_n3516# 7.7e-21
C1836 B7 a_636_n4294# 1.25417f
C1837 a_5288_n2434# a_5456_n2434# 2.18e-19
C1838 B0 a_11_46# 3.15e-19
C1839 a_3832_n2068# a_2995_n4294# 4.61e-19
C1840 A1 a_2254_n1194# 2.18e-20
C1841 a_894_n2068# B4 3.03e-19
C1842 a_3543_n2822# a_3368_n4255# 5.67e-19
C1843 a_541_n3308# a_n131_n1814# 2.21e-19
C1844 a_3795_n2734# a_3322_n4062# 0.010797f
C1845 a_798_n2434# a_1557_n2434# 0.031298f
C1846 A3 a_1261_n3080# 8.18e-21
C1847 a_2254_n2434# a_2422_n2434# 0.00792f
C1848 a_5773_n4294# a_4204_n3054# 1.52e-19
C1849 B1 a_143_n1036# 0.046267f
C1850 a_2350_n2068# B5 2.91e-19
C1851 a_5819_n2068# B8 0.033026f
C1852 Cin a_n131_n574# 0.001571f
C1853 a_4441_n3054# a_4204_n3054# 0.073551f
C1854 a_1968_n4294# a_2273_n2734# 0.14976f
C1855 a_2995_n4294# a_1647_n3054# 2.36e-19
C1856 DVDD a_1641_n3308# 0.160791f
C1857 a_5402_174# a_5456_46# 0.044963f
C1858 a_3874_n1220# B14 0.013754f
C1859 a_101_n3674# a_11_n3308# 0.006823f
C1860 DVDD a_541_n1194# 0.002071f
C1861 a_1201_n574# a_3543_n342# 3.23e-20
C1862 a_n131_n574# a_3669_n342# 6.1e-20
C1863 a_1201_n1814# a_2908_n600# 1.16e-19
C1864 a_636_n1814# a_n131_n1814# 0.044377f
C1865 A15 a_3765_n3080# 2.02e-21
C1866 a_4204_n3054# a_4000_n2068# 1.25e-20
C1867 a_4363_n3674# a_5402_n3546# 1.11e-20
C1868 a_143_n1036# a_1641_n828# 0.00341f
C1869 a_2273_n254# a_1467_n828# 1.07e-20
C1870 B3 a_n131_n1814# 0.00432f
C1871 a_2273_n2734# a_2459_n2734# 7.42e-19
C1872 B13 a_4691_n254# 0.002612f
C1873 a_3874_n1220# a_4363_46# 1.55e-21
C1874 B8 a_3765_n3080# 4.3e-20
C1875 A11 a_4691_n3974# 0.001028f
C1876 Cin a_3434_n1546# 1.05e-19
C1877 a_1647_n3054# a_1201_n4294# 1.02e-20
C1878 A0 a_147_n254# 0.001052f
C1879 a_143_n2276# a_1291_n3054# 8.48e-19
C1880 a_3226_n4062# a_2995_n4294# 0.101376f
C1881 a_1997_n3674# a_143_n3516# 4.76e-20
C1882 DVDD a_6153_46# 2.33e-19
C1883 B2 a_894_n1194# 7.33e-20
C1884 a_3946_174# a_4363_46# 0.06777f
C1885 a_2254_n1194# a_2315_n1775# 6.53e-19
C1886 a_798_n1194# a_636_n1814# 0.012687f
C1887 a_894_n828# a_101_n1194# 4.35e-21
C1888 a_1557_n1194# A3 0.791917f
C1889 A7 a_2422_n3308# 1.05e-19
C1890 a_3434_n1546# a_3669_n342# 0.055436f
C1891 a_3655_n1516# a_3543_n342# 0.011237f
C1892 a_143_n2276# a_541_n2434# 0.045338f
C1893 a_798_n1194# B3 2.55e-19
C1894 A4 a_n71_n3080# 0.081598f
C1895 DVDD a_1968_n1814# 0.307244f
C1896 B2 a_143_n1036# 0.662565f
C1897 B0 a_798_46# 0.078639f
C1898 Cin a_541_412# 0.088227f
C1899 S15 a_n131_n574# 3.89e-19
C1900 DVDD a_966_412# 7.01e-19
C1901 a_2273_n2734# a_2422_n2434# 2.27e-20
C1902 B14 a_6023_n1494# 0.002402f
C1903 A5 a_1641_n1194# 1.4e-21
C1904 B15 a_4363_n828# 0.020016f
C1905 a_2569_n4255# a_n131_n4294# 0.015565f
C1906 a_3543_n2822# a_6023_n2734# 6.93e-20
C1907 a_3543_n2822# a_3904_n3674# 0.008425f
C1908 DVDD a_6023_n574# 0.242051f
C1909 a_143_n2276# a_2569_n4255# 0.089244f
C1910 a_n131_n1814# a_2783_n1775# 8.19e-19
C1911 a_101_n2434# a_n131_n1814# 0.015023f
C1912 a_5855_n1814# a_3543_n342# 0.003681f
C1913 a_4691_n1814# a_3669_n342# 0.083702f
C1914 a_3874_n2460# B10 9.78e-20
C1915 A12 a_3765_n600# 4.94e-20
C1916 a_3874_20# a_4441_n1814# 9.91e-21
C1917 A8 a_5288_n2434# 5.43e-19
C1918 A3 a_1647_n574# 3.39e-19
C1919 a_3874_n2460# a_3434_n1546# 1.74e-20
C1920 A4 a_541_n3308# 3.08e-21
C1921 a_2273_n254# a_2350_412# 1.21e-20
C1922 a_1291_n1814# a_1201_n1814# 0.083702f
C1923 DVDD a_4523_n1814# 0.008551f
C1924 A7 a_2315_n4255# 0.002825f
C1925 a_315_n1814# a_636_n1814# 8e-20
C1926 B1 a_1641_n828# 9.06e-20
C1927 a_6023_n3974# B10 0.002402f
C1928 a_2995_n4294# a_3832_n2434# 8.24e-19
C1929 a_3946_n2306# a_4000_n2434# 0.046215f
C1930 a_3874_n2460# a_4363_n2434# 0.033252f
C1931 DVDD A13 0.443155f
C1932 a_185_n3308# a_541_n3308# 0.009846f
C1933 a_143_n2276# a_1997_n3674# 8.49e-20
C1934 A11 a_3832_n3674# 5.43e-19
C1935 a_3322_n1582# a_3226_n1582# 0.318695f
C1936 A12 a_5819_n1194# 1.17e-19
C1937 a_798_n1194# a_101_n2434# 9.75e-22
C1938 a_636_n3054# A3 0.00421f
C1939 a_143_n1036# a_1641_46# 8.74e-19
C1940 B5 a_2350_n2434# 7.33e-20
C1941 a_636_n1814# A4 4.8e-19
C1942 A5 A9 0.006192f
C1943 a_636_n3054# B9 2.79e-20
C1944 A9 a_4691_n2734# 9.63e-19
C1945 DVDD a_3685_n4255# 8.63e-19
C1946 a_2569_n3928# a_1968_n4294# 0.005193f
C1947 a_315_n4294# a_n71_n4320# 0.006406f
C1948 a_5819_n3674# a_3543_n2822# 0.001149f
C1949 B15 A14 2.69e-19
C1950 A15 B14 1.74e-19
C1951 a_4441_n3054# a_3669_n342# 4.02e-20
C1952 a_5773_n3054# a_3543_n342# 0.001891f
C1953 A7 a_1467_n3674# 5.03e-19
C1954 a_4204_n574# a_5192_n828# 2.69e-19
C1955 a_3543_n2822# a_2273_n2734# 3.18e-19
C1956 DVDD a_1467_n828# 4.94e-19
C1957 a_5819_n2068# a_2995_n4294# 0.091536f
C1958 a_5456_n2068# a_5402_n2306# 0.004108f
C1959 B6 a_315_n4294# 0.007771f
C1960 B14 a_5819_n828# 0.033026f
C1961 B14 B8 0.008756f
C1962 a_1557_n1194# a_1201_n574# 5.07e-20
C1963 a_636_n1814# a_1201_n1814# 0.105485f
C1964 a_101_n1194# a_636_n1814# 0.201352f
C1965 A15 a_4363_46# 1.4e-21
C1966 a_3543_n342# a_4363_n2068# 0.001068f
C1967 a_3946_n2306# a_3627_n2734# 3.01e-19
C1968 B3 a_1201_n1814# 0.081283f
C1969 a_2995_n4294# a_2543_n2734# 2.59e-19
C1970 a_5819_n2068# a_4204_n574# 1.77e-21
C1971 a_n41_n1814# B4 2.12e-19
C1972 B7 a_2254_n3674# 0.077341f
C1973 DVDD a_5402_174# 0.385125f
C1974 a_101_n1194# B3 7.19e-19
C1975 a_3655_n3996# a_2995_n4294# 0.042723f
C1976 a_101_46# a_n131_n574# 0.004436f
C1977 a_4204_n3054# a_5288_n2434# 1.66e-19
C1978 A7 B5 0.007762f
C1979 B7 A5 0.004004f
C1980 a_n131_n574# a_n71_n1840# 1.01e-20
C1981 a_1261_n600# a_1261_n1840# 0.002078f
C1982 a_3946_n2306# a_3861_n3080# 0.060379f
C1983 a_3874_n2460# a_4441_n3054# 0.01589f
C1984 a_2995_n4294# a_3765_n3080# 0.019426f
C1985 a_143_n2276# a_2497_n1775# 6.56e-19
C1986 A13 B13 1.25311f
C1987 a_5360_n1194# a_4697_n1194# 5.49e-20
C1988 a_1641_n2434# a_636_n3054# 0.033252f
C1989 a_1467_n2434# a_1557_n2434# 0.006958f
C1990 a_1997_n2434# a_101_n2434# 5.42e-21
C1991 a_5819_n3308# B8 5.74e-19
C1992 a_894_46# a_798_46# 0.005587f
C1993 a_101_n2434# A4 0.780011f
C1994 a_3874_n1220# a_3434_n1546# 1.72e-19
C1995 a_3946_n1066# a_3226_n1582# 4.55e-19
C1996 B1 a_1641_46# 0.019568f
C1997 a_6023_n3974# a_5773_n4294# 0.007234f
C1998 a_2422_n1194# a_2254_n1194# 0.00792f
C1999 a_1201_n1814# a_1291_n574# 2.26e-19
C2000 a_1201_n574# a_1647_n574# 0.001897f
C2001 a_1291_n4294# a_2995_n4294# 2.11e-19
C2002 a_3627_n254# a_3669_n342# 0.008516f
C2003 a_2543_n254# a_3765_n600# 1.71e-20
C2004 a_3874_n2460# a_4000_n2068# 0.112124f
C2005 a_3627_n2734# a_1201_n3054# 1.71e-20
C2006 a_3946_n2306# a_3904_n2434# 0.055111f
C2007 a_2543_n2734# a_1201_n4294# 0.008516f
C2008 DVDD a_2350_n2068# 4.94e-19
C2009 B12 a_3543_n342# 4.07e-19
C2010 a_185_n828# a_143_n1036# 0.091015f
C2011 DVDD a_2422_n3308# 6.64e-19
C2012 a_3946_174# a_3434_n1546# 2.72e-21
C2013 a_3946_n1066# a_4000_n2434# 6.4e-20
C2014 a_3434_n4026# a_n131_n4294# 1.44e-19
C2015 a_143_n2276# a_3434_n4026# 1.05e-19
C2016 a_3946_n3546# a_3904_n3674# 0.051953f
C2017 a_3874_n3700# a_4000_n3308# 0.112124f
C2018 a_3861_n3080# a_1201_n3054# 4.08e-20
C2019 a_3765_n3080# a_1201_n4294# 6.3e-20
C2020 a_3669_n2822# a_n131_n4294# 1.68e-20
C2021 B11 a_4691_n3054# 0.001447f
C2022 DVDD a_2350_412# 4.94e-19
C2023 B5 a_2273_n254# 0.002237f
C2024 Cin a_1641_412# 0.010774f
C2025 a_143_n2276# a_3669_n2822# 2.26e-20
C2026 a_143_n2276# a_1641_n1194# 0.001593f
C2027 B7 a_n71_n4320# 3.52e-21
C2028 DVDD a_n41_n3054# 0.244494f
C2029 DVDD a_4000_n3308# 0.154852f
C2030 a_3874_n1220# a_4691_n1814# 6.24e-19
C2031 a_3322_n1582# a_3904_n2434# 2.41e-19
C2032 a_101_n1194# a_101_n2434# 0.002006f
C2033 a_3226_n4062# a_3368_n4255# 0.005572f
C2034 a_5402_n2306# A9 1.36e-19
C2035 a_315_n4294# a_n131_n4294# 0.003681f
C2036 a_1291_n4294# a_1201_n4294# 0.083702f
C2037 B6 B7 0.003904f
C2038 B13 a_5402_174# 7.19e-19
C2039 A10 a_5819_n3308# 0.011602f
C2040 a_6023_n1814# A8 7.55e-19
C2041 a_541_n2068# a_143_n2276# 0.091602f
C2042 a_101_46# a_541_412# 0.004108f
C2043 a_4691_n3054# a_4204_n3054# 0.016475f
C2044 B7 a_143_n3516# 0.020606f
C2045 Cin a_n131_n1814# 0.524204f
C2046 a_1968_n4294# a_1557_n3674# 0.116264f
C2047 a_3322_n1582# a_3736_412# 4.54e-21
C2048 a_3226_n1582# a_3368_n1775# 0.005572f
C2049 B14 a_3861_n600# 7.86e-19
C2050 a_3736_n1194# a_4000_n1194# 8.12e-20
C2051 DVDD a_2315_n4255# 0.1905f
C2052 a_6023_n1814# a_5773_n1814# 0.025037f
C2053 a_6023_n3054# a_5773_n3054# 0.025037f
C2054 a_3736_n3674# a_3322_n4062# 4.57e-19
C2055 a_2908_n600# a_3543_n342# 0.06244f
C2056 B14 a_5360_46# 1.22e-20
C2057 B15 a_2254_n1194# 1.77e-20
C2058 a_2497_n1775# a_1968_n1814# 4.9e-19
C2059 a_143_n2276# A9 1.35e-19
C2060 a_5456_n3674# a_5402_n3546# 0.044963f
C2061 a_3832_n3308# a_4000_n3308# 2.18e-19
C2062 a_3946_n3546# a_2273_n2734# 8.35e-21
C2063 a_143_n2276# a_2363_n254# 9.97e-20
C2064 a_3946_n1066# a_3861_n3080# 2.93e-22
C2065 DVDD a_6153_n3674# 2.33e-19
C2066 Cin a_798_n1194# 1.17e-20
C2067 a_1641_n3674# a_1557_n3674# 0.06777f
C2068 a_4441_n574# a_2908_n600# 5.2e-21
C2069 DVDD a_3832_412# 4.94e-19
C2070 a_3669_n342# a_4697_n1194# 9.84e-21
C2071 a_3543_n342# a_5192_n1194# 1.65e-19
C2072 B14 a_2995_n4294# 7.21e-19
C2073 a_3946_n1066# a_3904_n2434# 1.25e-21
C2074 a_3874_20# a_3543_n342# 5.56e-19
C2075 B1 a_2422_46# 6.11e-20
C2076 B0 a_147_n1494# 2.47e-20
C2077 a_1641_n2068# a_636_n1814# 1.77e-21
C2078 a_5402_n2306# a_5402_n3546# 0.007891f
C2079 a_3543_n342# a_5456_n2434# 0.001136f
C2080 a_1641_n2068# B3 9.06e-20
C2081 S15 a_n131_n1814# 0.011587f
C2082 A15 a_3434_n1546# 0.00356f
C2083 B14 a_4204_n574# 0.662565f
C2084 B7 a_n131_n4294# 0.00432f
C2085 a_185_n2068# a_143_n1036# 1.77e-21
C2086 B7 a_143_n2276# 6.73e-19
C2087 B8 B10 0.013937f
C2088 a_3874_20# a_4441_n574# 0.01589f
C2089 DVDD B5 0.594006f
C2090 a_5819_n3308# a_2995_n4294# 1.77e-21
C2091 DVDD a_4000_n828# 0.154852f
C2092 a_5456_n3308# a_5402_n2306# 4.9e-19
C2093 a_147_n3974# B4 2.47e-20
C2094 B11 a_3322_n4062# 0.040998f
C2095 a_798_n2434# A2 2.18e-20
C2096 a_n131_n1814# a_n131_n3054# 0.001229f
C2097 a_4204_n574# a_4363_46# 8.74e-19
C2098 a_n41_n574# a_n71_n600# 0.025037f
C2099 DVDD a_n41_n574# 0.244494f
C2100 a_143_n2276# a_2350_n828# 3.53e-20
C2101 a_3946_n2306# B9 0.17279f
C2102 a_4691_n1814# A15 0.007493f
C2103 a_2273_n2734# a_1647_n3054# 3.8e-19
C2104 A2 a_541_n828# 0.011819f
C2105 B7 a_1641_n3308# 0.020016f
C2106 B2 a_185_n828# 0.033026f
C2107 a_3946_174# a_3627_n254# 3.01e-19
C2108 a_2995_n4294# a_4697_n2434# 1.77e-20
C2109 a_3874_n2460# a_5288_n2434# 2.34e-19
C2110 a_3946_n2306# a_5192_n2434# 3.2e-20
C2111 DVDD a_3368_n1448# 4.92e-19
C2112 a_3368_n3928# a_2995_n4294# 0.001315f
C2113 B13 a_3832_412# 2.91e-19
C2114 A13 a_3904_46# 0.114466f
C2115 a_3434_n4026# a_3685_n4255# 4.9e-19
C2116 a_966_n2434# a_143_n3516# 1.96e-19
C2117 a_5456_n2434# a_5819_n2434# 0.008475f
C2118 a_3669_n2822# a_3685_n4255# 2.79e-19
C2119 a_3543_n2822# a_4523_n4294# 0.002766f
C2120 a_3322_n4062# a_4204_n3054# 0.01799f
C2121 B9 a_3322_n1582# 0.002237f
C2122 A3 a_1201_n3054# 2.02e-21
C2123 a_1467_n2068# a_636_n3054# 7.45e-20
C2124 A10 B10 1.27934f
C2125 A7 a_3874_n3700# 2.02e-20
C2126 DVDD a_5456_46# 8.16e-19
C2127 Cin a_1201_n1814# 0.01502f
C2128 a_101_n3674# a_n131_n1814# 2.04e-19
C2129 a_5855_n3054# a_3543_n342# 2.76e-19
C2130 DVDD A7 0.470479f
C2131 a_1557_46# a_2254_46# 0.055111f
C2132 a_3543_n2822# a_1557_n3674# 1.19e-20
C2133 a_3226_n4062# a_2273_n2734# 2.95e-19
C2134 A6 a_147_n3974# 0.001052f
C2135 a_5402_n1066# B14 0.181244f
C2136 B5 a_1291_n3054# 0.05645f
C2137 DVDD a_966_n1194# 9.02e-20
C2138 a_5456_412# a_5819_412# 0.009846f
C2139 a_1201_n574# a_3765_n600# 0.001811f
C2140 a_n131_n574# a_3861_n600# 7.7e-20
C2141 A11 a_3946_n2306# 3.41e-19
C2142 a_3874_n1220# a_n131_n1814# 1.63e-21
C2143 a_1557_n1194# a_2908_n600# 6.6e-20
C2144 a_636_n1814# a_3543_n342# 1.63e-21
C2145 a_1467_n2434# a_2995_n4294# 3.6e-21
C2146 A15 a_4441_n3054# 8.18e-21
C2147 a_143_n1036# a_2254_n1194# 2.01e-19
C2148 a_2273_n254# a_1997_n828# 0.003825f
C2149 a_5773_n4294# B8 8.21e-21
C2150 a_966_n828# a_n131_n1814# 3.51e-20
C2151 DVDD a_2790_n3928# 4.92e-19
C2152 B3 a_3543_n342# 1.25e-20
C2153 a_11_n3674# a_101_n3674# 0.006958f
C2154 a_1291_n1814# a_1261_n3080# 9.75e-20
C2155 a_147_n254# a_1201_n574# 2.05e-20
C2156 DVDD a_2273_n254# 1.16079f
C2157 a_185_n2434# a_101_n2434# 0.067562f
C2158 A8 a_3543_n342# 0.012262f
C2159 a_101_46# a_n131_n1814# 2.69e-19
C2160 a_3874_n2460# a_4691_n3054# 0.006212f
C2161 a_143_n2276# a_2569_n1448# 3.99e-19
C2162 A15 a_4000_n2068# 8.69e-21
C2163 a_5288_n828# a_5360_n1194# 0.004869f
C2164 a_5288_n3674# B10 7.33e-20
C2165 a_n131_n1814# a_n71_n1840# 0.188784f
C2166 a_3946_n1066# a_4363_n1194# 0.06777f
C2167 a_3946_n1066# A3 2.18e-20
C2168 a_4441_n1814# a_3669_n342# 0.188936f
C2169 a_5773_n1814# a_3543_n342# 0.188784f
C2170 a_3655_n1516# a_3765_n600# 2.4e-19
C2171 a_3434_n1546# a_3861_n600# 5.85e-21
C2172 a_143_n2276# a_966_n2434# 4.46e-19
C2173 a_4363_n3674# B9 2.95e-21
C2174 A4 a_n131_n3054# 0.025968f
C2175 a_798_n1194# a_966_n828# 0.007578f
C2176 a_3946_n1066# B9 2.43e-20
C2177 A7 a_1291_n3054# 7.81e-20
C2178 A12 a_5288_46# 5.43e-19
C2179 B12 a_5192_46# 6.11e-20
C2180 S15 a_1201_n1814# 0.003272f
C2181 a_3655_n3996# a_3904_n3674# 6.53e-19
C2182 a_798_n1194# a_101_46# 1.16e-19
C2183 a_3861_n3080# a_4691_n2734# 9.28e-20
C2184 a_3765_n3080# a_6023_n2734# 2.05e-20
C2185 a_3669_n2822# a_4000_n3308# 4.28e-19
C2186 a_3765_n3080# a_3904_n3674# 4.56e-19
C2187 A3 a_1261_n1840# 0.084607f
C2188 a_3322_n1582# a_1201_n574# 2.76e-20
C2189 A10 a_5773_n4294# 0.081598f
C2190 a_3543_n342# a_2783_n1775# 3.15e-20
C2191 a_6023_n1814# a_3669_n342# 2.66e-19
C2192 a_1557_n2434# a_n131_n1814# 0.001955f
C2193 B2 a_185_n2068# 5.74e-19
C2194 a_3946_174# a_3832_46# 3.53e-19
C2195 a_3874_20# a_4000_46# 0.045338f
C2196 a_1201_n1814# a_n131_n3054# 5.47e-21
C2197 a_143_n2276# a_1261_n600# 0.001345f
C2198 A8 a_5819_n2434# 0.050725f
C2199 a_3874_n2460# a_4441_n1814# 5.78e-19
C2200 a_2995_n4294# a_3434_n1546# 0.011854f
C2201 a_541_n3308# a_798_n3674# 0.02283f
C2202 a_3946_n2306# a_3655_n1516# 9.88e-20
C2203 A5 a_3904_n2434# 9.68e-20
C2204 A11 a_636_n4294# 2.02e-20
C2205 a_1641_n2434# a_636_n4294# 1.55e-21
C2206 B3 a_1261_n3080# 3.66e-21
C2207 a_5402_n2306# a_4000_n2434# 5.42e-21
C2208 a_2995_n4294# a_4363_n2434# 0.005715f
C2209 A4 a_101_n3674# 6.66e-20
C2210 a_1968_n4294# a_3543_n2822# 1.44e-19
C2211 A3 a_2254_46# 1.29e-20
C2212 A11 a_4363_n3674# 0.051667f
C2213 A1 a_n131_n574# 0.022989f
C2214 a_4204_n574# a_3434_n1546# 8.25e-20
C2215 a_3322_n1582# a_3655_n1516# 0.236061f
C2216 a_3874_n3700# a_4691_n4294# 6.24e-19
C2217 a_5402_174# a_5819_46# 0.067562f
C2218 a_4691_n1814# a_2995_n4294# 0.006854f
C2219 a_4204_n3054# a_3543_n342# 1.24e-19
C2220 a_101_n3674# a_185_n3308# 0.030161f
C2221 a_2273_n2734# a_2543_n2734# 7.04e-19
C2222 a_2569_n1448# a_1968_n1814# 0.005193f
C2223 a_315_n1814# a_n71_n1840# 0.006406f
C2224 DVDD a_4691_n4294# 0.259723f
C2225 A9 a_4000_n3308# 8.69e-21
C2226 a_2790_n3928# a_2569_n4255# 0.007833f
C2227 a_143_n2276# a_3226_n1582# 0.00672f
C2228 a_1291_n4294# a_1261_n4320# 0.025037f
C2229 a_3655_n3996# a_2273_n2734# 2.02e-20
C2230 a_1557_n3674# a_3946_n3546# 0.001288f
C2231 B15 a_3765_n3080# 5.62e-22
C2232 A7 a_1997_n3674# 0.046632f
C2233 a_3765_n3080# a_2273_n2734# 3.67e-20
C2234 DVDD a_1997_n828# 0.154852f
C2235 a_6153_n2068# a_5402_n2306# 0.006823f
C2236 a_4691_n1814# a_4204_n574# 1.59e-20
C2237 A15 a_n131_n1814# 1.12e-19
C2238 DVDD a_3874_n3700# 1.042f
C2239 B11 a_4691_n3974# 0.002951f
C2240 A4 a_n71_n1840# 0.001911f
C2241 a_5360_n1194# a_3543_n342# 0.001991f
C2242 a_3874_n1220# a_1201_n1814# 1.36e-21
C2243 B0 a_147_n254# 0.002402f
C2244 a_1479_n254# a_1261_n600# 0.007234f
C2245 DVDD a_n71_n600# 0.176878f
C2246 a_3832_412# a_3904_46# 0.004869f
C2247 B4 a_n71_n3080# 0.226175f
C2248 a_636_n1814# a_1557_n1194# 0.287345f
C2249 a_636_n3054# a_n71_n3080# 0.063303f
C2250 a_101_n2434# a_1261_n3080# 0.005909f
C2251 a_1291_n4294# a_2273_n2734# 1.57e-19
C2252 a_3543_n342# a_5192_n2068# 4.28e-20
C2253 A8 a_6023_n3054# 0.007489f
C2254 a_3874_20# a_5192_46# 3.15e-19
C2255 a_3946_174# a_4697_46# 0.006958f
C2256 a_3946_n2306# a_3795_n2734# 6.28e-19
C2257 a_3874_n2460# a_3322_n4062# 3.49e-19
C2258 a_2995_n4294# a_3711_n2734# 9.55e-19
C2259 a_1557_n1194# B3 0.175017f
C2260 B7 a_2422_n3308# 3.18e-19
C2261 a_894_n2068# a_143_n3516# 3.3e-20
C2262 A15 a_4697_n1194# 5.03e-19
C2263 a_4204_n3054# a_5819_n2434# 1.55e-21
C2264 a_2995_n4294# a_4441_n3054# 0.004963f
C2265 a_101_n1194# a_101_46# 0.007891f
C2266 a_5402_n2306# a_3861_n3080# 0.004436f
C2267 a_n131_n574# a_2315_n1775# 5.6e-20
C2268 a_1201_n1814# a_n71_n1840# 3.93e-19
C2269 a_1201_n574# a_1261_n1840# 7.34e-21
C2270 a_5360_n1194# a_5288_n1194# 0.005587f
C2271 a_101_n1194# a_n71_n1840# 0.003994f
C2272 a_1997_n2434# a_1557_n2434# 0.046215f
C2273 A0 a_966_412# 1.05e-19
C2274 Cin a_798_46# 0.087504f
C2275 A2 a_n131_n574# 2.3e-19
C2276 DVDD a_1467_412# 5e-19
C2277 B0 a_894_412# 3.03e-19
C2278 a_101_n2434# a_798_n3674# 1.16e-19
C2279 a_1557_n2434# A4 0.001406f
C2280 B5 a_1641_n1194# 3.27e-20
C2281 a_5402_n1066# a_3434_n1546# 4.58e-20
C2282 a_3874_n1220# a_4441_n1814# 0.015611f
C2283 a_3946_n1066# a_3655_n1516# 0.027489f
C2284 a_3832_n3308# a_3874_n3700# 1.35e-20
C2285 a_3874_n2460# a_4697_n2068# 7.45e-20
C2286 a_3795_n254# a_3669_n342# 1.46e-22
C2287 a_2995_n4294# a_4000_n2068# 0.015774f
C2288 a_3946_n2306# a_4363_n2068# 0.030161f
C2289 a_3322_n4062# a_n131_n3054# 1.64e-19
C2290 a_3711_n254# a_3765_n600# 0.009339f
C2291 B12 a_3765_n600# 4.3e-20
C2292 DVDD a_3736_n2068# 6.64e-19
C2293 DVDD a_3832_n3308# 4.94e-19
C2294 DVDD a_4000_n1194# 8.16e-19
C2295 B8 a_5288_n2434# 7.33e-20
C2296 A6 a_n71_n3080# 0.001913f
C2297 a_3874_n3700# a_4697_n3308# 7.45e-20
C2298 a_3946_n3546# a_4363_n3308# 0.030161f
C2299 a_2273_n254# a_2422_412# 4.54e-21
C2300 a_3861_n3080# a_n131_n4294# 8.62e-20
C2301 a_1201_n574# a_2254_46# 4.74e-19
C2302 a_3226_n1582# a_1968_n1814# 3.07e-19
C2303 a_5360_n2434# A14 2.18e-20
C2304 a_143_n2276# a_3861_n3080# 3.22e-20
C2305 a_1997_n2068# A3 8.69e-21
C2306 a_1557_n2434# a_1201_n1814# 5.83e-20
C2307 B7 a_2315_n4255# 2.1e-19
C2308 DVDD a_1291_n3054# 0.238543f
C2309 a_636_n1814# B4 1.83e-19
C2310 DVDD a_4697_n3308# 4.94e-19
C2311 a_2350_n1194# A3 5.43e-19
C2312 a_3874_n1220# a_6023_n1814# 1.77e-19
C2313 a_636_n1814# a_636_n3054# 0.001068f
C2314 DVDD B13 0.565562f
C2315 A12 a_6153_46# 4.78e-19
C2316 B11 a_3832_n3674# 7.33e-20
C2317 A3 A5 0.001672f
C2318 a_636_n3054# B3 1.13e-19
C2319 a_1647_n4294# a_n131_n4294# 0.002766f
C2320 DVDD a_541_n2434# 8.16e-19
C2321 a_143_n2276# a_3904_n2434# 1.26e-19
C2322 A5 B9 2.72e-20
C2323 B5 A9 2.72e-20
C2324 A6 a_541_n3308# 0.011819f
C2325 A7 a_3669_n2822# 7.21e-20
C2326 a_2497_n1775# a_2273_n254# 0.005265f
C2327 B9 a_4691_n2734# 0.002612f
C2328 a_894_n2068# a_143_n2276# 5.19e-19
C2329 Cin a_3543_n342# 1.28e-19
C2330 a_6023_n3054# a_4204_n3054# 0.002038f
C2331 B15 B14 0.003904f
C2332 a_3434_n1546# a_3685_n1775# 4.9e-19
C2333 B7 a_1467_n3674# 6.45e-19
C2334 DVDD a_2569_n4255# 0.105346f
C2335 a_143_n2276# a_1557_46# 9.58e-19
C2336 a_4000_n3674# a_3322_n4062# 0.001323f
C2337 a_3322_n1582# a_3711_n254# 7.42e-19
C2338 a_3543_n342# a_3669_n342# 1.11131f
C2339 a_n131_n1814# a_3861_n600# 8.62e-20
C2340 a_2790_n3928# a_3434_n4026# 8.12e-20
C2341 a_2908_n600# a_3765_n600# 5.75e-19
C2342 A12 a_6023_n574# 0.007489f
C2343 a_6153_n3674# a_5402_n3546# 0.006958f
C2344 DVDD a_185_46# 0.003788f
C2345 B15 a_4363_46# 3.27e-20
C2346 a_143_n2276# a_2543_n254# 6.51e-20
C2347 a_101_46# a_11_46# 0.006958f
C2348 A15 a_1201_n1814# 7.21e-20
C2349 DVDD a_11_412# 5.28e-19
C2350 A11 a_2254_n3674# 9.68e-20
C2351 a_101_n2434# B4 0.181244f
C2352 a_101_n2434# a_636_n3054# 0.172114f
C2353 a_5773_n574# a_3543_n342# 0.001041f
C2354 a_4441_n574# a_3669_n342# 3.76e-19
C2355 a_636_n574# a_n131_n574# 0.289331f
C2356 a_3543_n342# a_5456_n1194# 0.001186f
C2357 DVDD a_1997_n3674# 8.16e-19
C2358 B7 B5 0.005115f
C2359 a_1641_n2434# A5 0.051667f
C2360 A13 A12 0.019542f
C2361 a_3874_20# a_3765_n600# 0.104793f
C2362 a_3874_n2460# a_3543_n342# 0.001496f
C2363 a_3946_n2306# a_2908_n600# 9.75e-22
C2364 a_966_46# a_798_46# 0.00792f
C2365 a_798_n2434# a_143_n1036# 1.17e-20
C2366 a_3543_n342# a_6153_n2434# 1.2e-19
C2367 S15 a_3543_n342# 3.74e-19
C2368 a_2254_n2434# a_n131_n574# 3.7e-21
C2369 A15 a_4441_n1814# 0.084607f
C2370 a_541_n828# a_143_n1036# 0.087066f
C2371 a_5288_n1194# a_5456_n1194# 2.18e-19
C2372 a_1997_n1194# a_1201_n1814# 0.001261f
C2373 a_2254_n3674# a_2350_n3674# 0.005587f
C2374 a_1997_n1194# a_101_n1194# 5.42e-21
C2375 a_3322_n1582# a_2908_n600# 0.024829f
C2376 Cin a_1997_412# 0.009966f
C2377 A1 a_1641_412# 0.011562f
C2378 DVDD a_2422_412# 6.64e-19
C2379 a_5456_46# a_5819_46# 0.008475f
C2380 a_2995_n4294# a_4697_n1194# 8.81e-21
C2381 DVDD a_4697_n828# 4.94e-19
C2382 A6 a_101_n2434# 0.003407f
C2383 a_n131_n1814# a_1201_n4294# 1.08e-20
C2384 a_2363_n254# a_2273_n254# 0.010797f
C2385 a_1647_n1814# a_n131_n1814# 0.002766f
C2386 a_147_n2734# a_n71_n3080# 0.007234f
C2387 A7 B7 1.25275f
C2388 a_5402_n2306# B9 7.19e-19
C2389 a_1557_46# a_1968_n1814# 2.72e-21
C2390 a_3946_174# a_3795_n254# 6.28e-19
C2391 a_5402_n2306# a_5192_n2434# 3.46e-19
C2392 A12 a_5402_174# 0.780011f
C2393 a_2995_n4294# a_5288_n2434# 4.74e-19
C2394 a_1968_n4294# a_3226_n4062# 3.07e-19
C2395 a_2497_n4255# a_2995_n4294# 9.03e-20
C2396 a_6023_n1814# B8 2.12e-19
C2397 DVDD a_5456_n2068# 0.1561f
C2398 DVDD a_2497_n1775# 8.63e-19
C2399 a_101_46# a_798_46# 0.057793f
C2400 a_3874_20# a_3322_n1582# 3.49e-19
C2401 A1 a_n131_n1814# 1.84e-20
C2402 a_1641_n2434# a_143_n3516# 8.74e-19
C2403 a_1641_n2068# a_1557_n2434# 0.030161f
C2404 a_3669_n2822# a_4691_n4294# 0.083702f
C2405 a_3543_n2822# a_5855_n4294# 0.003681f
C2406 a_3434_n1546# a_3904_n3674# 4.29e-21
C2407 a_143_n2276# A3 0.020847f
C2408 a_185_n1194# a_n131_n1814# 0.001149f
C2409 a_3434_n4026# a_3874_n3700# 1.72e-19
C2410 B7 a_2273_n254# 7.09e-22
C2411 Cin a_1557_n1194# 9.04e-19
C2412 a_143_n2276# B9 1.52e-20
C2413 a_3543_n2822# a_3946_n3546# 0.002594f
C2414 a_3669_n2822# a_3874_n3700# 0.105485f
C2415 DVDD a_3434_n4026# 0.301739f
C2416 DVDD a_3669_n2822# 0.365978f
C2417 a_2497_n4255# a_1201_n4294# 2.79e-19
C2418 A13 a_1557_46# 2.18e-20
C2419 DVDD a_1641_n1194# 0.001386f
C2420 a_1201_n1814# a_3861_n600# 6.1e-20
C2421 a_1557_n1194# a_3669_n342# 9.92e-21
C2422 a_3946_n1066# a_2908_n600# 0.052161f
C2423 a_3874_n1220# a_3543_n342# 0.044242f
C2424 a_1997_n2434# a_2995_n4294# 8.26e-19
C2425 A13 a_3736_412# 1.05e-19
C2426 a_4697_46# a_5360_46# 5.49e-20
C2427 a_4204_n3054# a_5288_n2068# 3.3e-20
C2428 DVDD a_3904_46# 0.247054f
C2429 a_5360_n3674# a_3543_n2822# 0.001991f
C2430 a_2273_n254# a_2350_n828# 2.27e-19
C2431 DVDD a_315_n4294# 0.009643f
C2432 a_n71_n3080# a_1201_n3054# 2.84e-19
C2433 a_1261_n3080# a_n131_n3054# 0.041433f
C2434 a_3946_174# a_3543_n342# 7.63e-19
C2435 a_2995_n4294# a_4691_n3054# 0.001398f
C2436 a_3874_n2460# a_6023_n3054# 4.33e-19
C2437 a_541_n2068# DVDD 0.1561f
C2438 a_143_n2276# a_n41_n1814# 7.37e-19
C2439 a_3874_n1220# a_4441_n574# 5.78e-19
C2440 a_5819_n3674# B10 0.021045f
C2441 a_5360_n1194# a_5456_n828# 0.02283f
C2442 a_n131_n1814# a_2315_n1775# 0.011237f
C2443 a_3946_n1066# a_5192_n1194# 3.2e-20
C2444 a_3874_n1220# a_5288_n1194# 2.34e-19
C2445 B15 a_3434_n1546# 0.002893f
C2446 A2 a_n131_n1814# 0.02685f
C2447 A11 a_n131_n4294# 1.12e-19
C2448 A11 a_143_n2276# 1.35e-19
C2449 a_4441_n1814# a_3861_n600# 9.27e-21
C2450 A9 a_3874_n3700# 0.004204f
C2451 a_3946_174# a_4441_n574# 0.002379f
C2452 a_2422_n3674# a_2995_n4294# 1.79e-19
C2453 a_143_n2276# a_1641_n2434# 0.004093f
C2454 a_3832_n3308# a_3669_n2822# 1.5e-20
C2455 DVDD A9 0.460573f
C2456 B15 a_4363_n2434# 2.95e-21
C2457 A10 a_3322_n4062# 5.21e-20
C2458 a_798_n2434# B2 1.17e-20
C2459 a_4204_n574# a_4697_46# 9.38e-21
C2460 a_3543_n2822# a_5192_n3308# 3.51e-20
C2461 A3 a_1968_n1814# 0.00356f
C2462 a_315_n574# a_n71_n600# 0.006406f
C2463 DVDD a_315_n574# 0.006628f
C2464 A0 a_n41_n574# 0.007489f
C2465 a_3946_n2306# A8 0.001406f
C2466 a_636_n1814# a_3322_n1582# 1.14e-21
C2467 a_4691_n1814# B15 0.056553f
C2468 a_3669_n342# a_4691_n1494# 0.002666f
C2469 a_3543_n342# a_6023_n1494# 0.002687f
C2470 B2 a_541_n828# 0.017703f
C2471 a_4441_n574# a_4523_n574# 0.006406f
C2472 A2 a_798_n1194# 0.114467f
C2473 a_1201_n1814# a_1201_n4294# 2.45e-20
C2474 a_541_n3308# a_966_n3308# 1.31e-19
C2475 a_2422_n3674# a_1201_n4294# 5.8e-19
C2476 a_1647_n1814# a_1201_n1814# 0.002223f
C2477 a_2995_n4294# a_4441_n1814# 0.009494f
C2478 a_798_n3674# a_894_n3308# 0.004869f
C2479 a_143_n2276# a_1201_n574# 0.002526f
C2480 a_1557_n1194# a_n131_n3054# 2.93e-22
C2481 A13 a_4000_412# 0.011819f
C2482 B13 a_3904_46# 0.077428f
C2483 a_143_n2276# a_2350_n3674# 1.03e-20
C2484 a_3874_20# a_4691_n574# 0.006212f
C2485 B3 a_1201_n3054# 5.62e-22
C2486 a_2569_n4255# a_3434_n4026# 3.07e-19
C2487 B7 a_3874_n3700# 2.79e-20
C2488 a_101_n3674# a_798_n3674# 0.057934f
C2489 a_n71_n4320# a_147_n3974# 0.007234f
C2490 DVDD a_5819_46# 0.001386f
C2491 a_3736_n2068# A9 1.05e-19
C2492 A1 a_1201_n1814# 0.001673f
C2493 a_3226_n4062# a_3543_n2822# 0.015332f
C2494 a_4000_n1194# A9 6.84e-21
C2495 a_4204_n574# a_4441_n1814# 5.74e-19
C2496 DVDD B7 0.610447f
C2497 a_1557_46# a_2350_412# 4.35e-21
C2498 a_3874_20# a_2254_46# 2.15e-20
C2499 B6 a_147_n3974# 0.002402f
C2500 a_3874_n3700# a_6023_n4294# 1.77e-19
C2501 a_5192_n3674# a_4204_n3054# 1.32e-19
C2502 a_636_n3054# a_3874_n2460# 0.001289f
C2503 a_6023_n1814# a_2995_n4294# 7.37e-19
C2504 a_636_n574# a_1641_412# 0.12395f
C2505 a_1291_n1814# a_1261_n1840# 0.025037f
C2506 a_2790_n1448# a_2569_n1775# 0.007833f
C2507 DVDD a_6023_n4294# 0.263648f
C2508 a_1997_n828# a_2350_n828# 2.18e-19
C2509 a_143_n2276# a_3655_n1516# 6.51e-19
C2510 a_3368_n1448# a_3226_n1582# 0.007833f
C2511 a_3177_n1814# a_3434_n1546# 2.84e-19
C2512 B11 a_3946_n2306# 4.05e-20
C2513 a_101_n1194# a_185_n1194# 0.067562f
C2514 a_3874_n3700# a_5402_n3546# 0.201352f
C2515 B15 a_4441_n3054# 3.66e-21
C2516 a_3765_n3080# a_2459_n2734# 9.58e-21
C2517 DVDD a_2350_n828# 4.94e-19
C2518 A15 a_3543_n342# 0.004783f
C2519 DVDD a_5402_n3546# 0.382636f
C2520 a_6023_n1814# a_4204_n574# 1.35e-19
C2521 a_185_n3674# a_101_n3674# 0.067562f
C2522 a_3832_n3674# a_4000_n3674# 2.18e-19
C2523 a_5819_n828# a_3543_n342# 5.74e-19
C2524 a_11_n1194# a_n131_n1814# 1.33e-19
C2525 a_636_n574# a_n131_n1814# 5.56e-19
C2526 B11 a_3322_n1582# 7.09e-22
C2527 a_1479_n254# a_1201_n574# 0.004527f
C2528 a_2273_n254# a_1261_n600# 6.57e-19
C2529 a_143_n1036# a_n131_n574# 0.182595f
C2530 B8 a_3543_n342# 0.015549f
C2531 B4 a_n131_n3054# 0.059236f
C2532 A2 A4 0.00475f
C2533 a_1557_n2434# a_1261_n3080# 0.002379f
C2534 a_636_n3054# a_n131_n3054# 0.289331f
C2535 a_101_n2434# a_1201_n3054# 0.003561f
C2536 a_5360_n3674# a_3946_n3546# 0.031298f
C2537 a_3946_n2306# a_4204_n3054# 0.057421f
C2538 a_2995_n4294# a_3322_n4062# 0.072877f
C2539 a_3946_n1066# B3 2.32e-20
C2540 DVDD a_5456_n3308# 0.1561f
C2541 A15 a_4441_n574# 1.75e-19
C2542 a_1479_n3974# a_2995_n4294# 1.33e-19
C2543 a_1201_n1814# a_2315_n1775# 0.024621f
C2544 a_5402_n2306# a_5773_n3054# 0.003994f
C2545 a_1201_n574# a_1968_n1814# 1.81e-21
C2546 A12 a_5456_46# 0.047225f
C2547 B7 a_1291_n3054# 0.001447f
C2548 B12 a_5288_46# 7.33e-20
C2549 a_636_n1814# a_1261_n1840# 0.015611f
C2550 a_2254_n2434# a_n131_n1814# 0.002327f
C2551 A2 a_1201_n1814# 1.6e-19
C2552 a_11_n828# a_n131_n1814# 9e-21
C2553 A2 a_101_n1194# 0.780011f
C2554 A14 a_5192_n828# 1.05e-19
C2555 a_5402_n1066# a_4441_n1814# 0.005934f
C2556 B3 a_1261_n1840# 0.2191f
C2557 a_3226_n1582# a_2273_n254# 3.13e-19
C2558 a_2995_n4294# a_4697_n2068# 8.12e-20
C2559 a_3322_n4062# a_1201_n4294# 7.77e-20
C2560 B4 a_101_n3674# 6.9e-19
C2561 a_636_n3054# a_101_n3674# 1.11e-19
C2562 a_3946_174# a_4000_46# 0.046215f
C2563 a_1641_n2068# a_2995_n4294# 3.36e-19
C2564 B8 a_5819_n2434# 0.021045f
C2565 A10 a_3543_n342# 8.62e-20
C2566 a_1479_n3974# a_1201_n4294# 0.002666f
C2567 a_147_n3974# a_n131_n4294# 0.002687f
C2568 A6 a_n131_n3054# 2.3e-19
C2569 B5 a_3904_n2434# 1.77e-20
C2570 B11 a_636_n4294# 2.79e-20
C2571 a_4204_n574# a_5288_n828# 2.9e-19
C2572 a_3322_n1582# a_5360_n1194# 2.74e-19
C2573 a_147_n1494# a_n71_n1840# 0.007234f
C2574 a_5819_n2068# A14 6.72e-19
C2575 a_3434_n1546# a_2569_n1775# 3.07e-19
C2576 a_185_n828# a_541_n828# 0.009846f
C2577 DVDD a_5288_n3308# 4.94e-19
C2578 DVDD a_2569_n1448# 2.55e-19
C2579 a_1557_n1194# a_1557_n2434# 0.0016f
C2580 a_1291_n574# a_1261_n1840# 9.75e-20
C2581 B11 a_4363_n3674# 0.019568f
C2582 B1 a_n131_n574# 0.033034f
C2583 a_5360_n3674# a_5192_n3308# 0.007578f
C2584 A9 a_3736_n2434# 7.66e-19
C2585 a_1467_n2068# a_143_n2276# 9.76e-20
C2586 B4 a_n71_n1840# 0.001358f
C2587 a_3226_n4062# a_3946_n3546# 4.55e-19
C2588 Cin a_3765_n600# 1.95e-20
C2589 a_3655_n3996# a_3543_n2822# 0.011237f
C2590 a_3434_n4026# a_3669_n2822# 0.055436f
C2591 a_3543_n2822# a_3765_n3080# 6.83e-19
C2592 A6 a_101_n3674# 0.780011f
C2593 B7 a_1997_n3674# 0.005557f
C2594 A10 a_5819_n2434# 4.33e-21
C2595 B15 a_n131_n1814# 1.25e-20
C2596 a_4363_n3674# a_4204_n3054# 9.15e-19
C2597 a_3669_n342# a_3765_n600# 0.15552f
C2598 a_3543_n342# a_3861_n600# 0.001745f
C2599 DVDD a_1261_n600# 0.173165f
C2600 A0 a_n71_n600# 0.081598f
C2601 DVDD A0 0.47691f
C2602 A5 a_n71_n3080# 1.38e-21
C2603 a_3832_412# a_4000_412# 2.18e-19
C2604 B8 a_6023_n3054# 0.056561f
C2605 a_3946_174# a_5192_46# 3.2e-20
C2606 a_3874_20# a_5288_46# 2.34e-19
C2607 a_1291_n1814# A5 7.81e-20
C2608 a_1557_n1194# A15 2.18e-20
C2609 a_2254_n2434# a_1997_n2434# 0.023012f
C2610 a_1557_n2434# B4 3.07e-19
C2611 a_4441_n574# a_3861_n600# 0.041433f
C2612 a_636_n3054# a_1557_n2434# 0.287408f
C2613 a_5773_n574# a_3765_n600# 2.84e-19
C2614 B15 a_4697_n1194# 6.45e-19
C2615 a_636_n574# a_1201_n1814# 7.1e-20
C2616 a_3946_n1066# a_5360_n1194# 0.031298f
C2617 a_5402_n1066# a_5288_n828# 4.35e-21
C2618 a_101_n1194# a_11_n1194# 0.006958f
C2619 a_101_n1194# a_636_n574# 1.11e-19
C2620 a_3368_n3928# a_1968_n4294# 8.12e-20
C2621 A11 a_4000_n3308# 0.011819f
C2622 Cin a_894_412# 2.96e-19
C2623 B2 a_n131_n574# 7.86e-19
C2624 A1 a_798_46# 0.001236f
C2625 B0 a_966_412# 3.18e-19
C2626 a_3946_n2306# a_3669_n342# 5.83e-20
C2627 a_2995_n4294# a_3543_n342# 0.330594f
C2628 a_11_n2068# a_n131_n1814# 3.89e-20
C2629 A9 a_3669_n2822# 0.001673f
C2630 DVDD a_3226_n1582# 0.108834f
C2631 Cin a_3322_n1582# 9.39e-19
C2632 a_n71_n4320# a_n71_n3080# 0.001197f
C2633 a_3736_n828# a_2908_n600# 0.007696f
C2634 A15 a_4000_46# 6.84e-21
C2635 a_541_n2434# a_966_n2434# 8.12e-20
C2636 S15 a_3765_n600# 9.75e-20
C2637 a_2422_n1194# a_1201_n1814# 5.8e-19
C2638 a_5456_n1194# a_5819_n1194# 0.008475f
C2639 a_2497_n4255# a_2273_n2734# 0.005265f
C2640 a_1997_n1194# a_1557_n1194# 0.046215f
C2641 a_1557_46# a_2273_n254# 0.008526f
C2642 a_11_n828# a_101_n1194# 0.006823f
C2643 DVDD a_4000_n2434# 8.16e-19
C2644 B6 a_n71_n3080# 0.001373f
C2645 a_4204_n574# a_3543_n342# 0.012648f
C2646 a_3322_n1582# a_3669_n342# 0.471487f
C2647 a_2995_n4294# a_4441_n574# 4.2e-19
C2648 A10 a_6023_n3054# 7.55e-19
C2649 a_5360_n2434# B14 1.17e-20
C2650 a_2350_n1194# B3 7.33e-20
C2651 a_143_n2276# a_2908_n600# 0.001132f
C2652 a_143_n3516# a_n71_n3080# 0.001762f
C2653 a_147_n2734# a_n131_n3054# 0.002789f
C2654 a_2543_n254# a_2273_n254# 7.04e-19
C2655 a_1479_n2734# a_1261_n3080# 0.007234f
C2656 a_3177_n1814# a_n131_n1814# 8.29e-19
C2657 a_3874_n2460# a_3946_n2306# 0.287408f
C2658 B12 a_6153_46# 3.15e-19
C2659 DVDD A12 0.460364f
C2660 A15 a_4691_n1494# 0.001028f
C2661 A3 B5 0.00374f
C2662 B3 A5 0.007762f
C2663 a_4204_n574# a_4441_n574# 0.073551f
C2664 a_5402_n2306# a_5456_n2434# 0.044963f
C2665 a_3322_n4062# a_3368_n4255# 0.006879f
C2666 a_2995_n4294# a_5819_n2434# 0.033252f
C2667 a_4204_n574# a_5288_n1194# 1.28e-19
C2668 B6 a_541_n3308# 0.017703f
C2669 B5 B9 0.001479f
C2670 B7 a_3669_n2822# 1.03e-20
C2671 DVDD a_6153_n2068# 5.28e-19
C2672 a_4691_n3974# a_2995_n4294# 5.95e-20
C2673 a_4441_n4294# a_4691_n4294# 0.025037f
C2674 A14 B14 1.27934f
C2675 a_3669_n2822# a_6023_n4294# 2.66e-19
C2676 a_143_n3516# a_541_n3308# 0.087066f
C2677 a_143_n1036# a_1641_412# 1.97e-19
C2678 A2 a_798_46# 1.29e-20
C2679 a_2995_n4294# a_1261_n3080# 7.81e-19
C2680 a_894_n1194# a_n131_n1814# 1.41e-19
C2681 a_3655_n3996# a_3946_n3546# 0.027489f
C2682 a_3434_n4026# a_5402_n3546# 4.58e-20
C2683 a_4441_n4294# a_3874_n3700# 0.015611f
C2684 S15 a_3322_n1582# 7.55e-19
C2685 DVDD a_3627_n2734# 2.46e-19
C2686 a_541_n3674# a_798_n3674# 0.023012f
C2687 B12 a_6023_n574# 0.056561f
C2688 Cin a_3946_n1066# 1.42e-20
C2689 a_3765_n3080# a_3946_n3546# 5.07e-20
C2690 a_3861_n3080# a_3874_n3700# 0.003854f
C2691 a_3669_n2822# a_5402_n3546# 0.003559f
C2692 DVDD a_4441_n4294# 0.183885f
C2693 A2 a_185_n2434# 1.15e-19
C2694 DVDD a_541_46# 0.002071f
C2695 A0 a_185_46# 0.050725f
C2696 a_5360_n2434# a_4697_n2434# 5.49e-20
C2697 B15 a_1201_n1814# 1.03e-20
C2698 DVDD a_3861_n3080# 1.67598f
C2699 a_2783_n4255# a_n131_n4294# 8.19e-19
C2700 B11 a_2254_n3674# 1.77e-20
C2701 a_143_n2276# a_2783_n4255# 1.1e-19
C2702 A0 a_11_412# 5.12e-20
C2703 a_101_n2434# A5 1.36e-19
C2704 a_3946_n1066# a_3669_n342# 0.044539f
C2705 a_3874_n1220# a_3765_n600# 1.04e-19
C2706 a_5402_n1066# a_3543_n342# 0.034089f
C2707 a_2422_n3674# a_2273_n2734# 4.57e-19
C2708 a_143_n1036# a_n131_n1814# 0.012648f
C2709 a_5819_n3308# a_3543_n2822# 5.74e-19
C2710 A4 a_11_n2068# 5.12e-20
C2711 a_798_n1194# a_894_n1194# 0.005587f
C2712 Cin a_1261_n1840# 1.44e-20
C2713 a_n71_n3080# a_n131_n4294# 0.001041f
C2714 a_1641_n2434# B5 0.019568f
C2715 a_1261_n3080# a_1201_n4294# 3.76e-19
C2716 a_n131_n3054# a_1201_n3054# 0.197466f
C2717 A13 B12 1.74e-19
C2718 DVDD a_1647_n4294# 0.008551f
C2719 B13 A12 2.69e-19
C2720 a_143_n2276# a_n71_n3080# 1.52e-19
C2721 a_3946_174# a_3765_n600# 0.076462f
C2722 DVDD a_3904_n2434# 0.247054f
C2723 a_1467_46# a_798_46# 5.49e-20
C2724 a_185_n3674# a_541_n3674# 0.008475f
C2725 a_2995_n4294# a_6023_n3054# 1.35e-19
C2726 a_894_n2068# DVDD 4.94e-19
C2727 a_143_n2276# a_1291_n1814# 0.011866f
C2728 a_5456_n828# a_5819_n828# 0.009846f
C2729 a_1557_46# a_1997_n828# 5.56e-19
C2730 a_n131_n1814# a_2569_n1775# 0.015565f
C2731 a_5402_n1066# a_5288_n1194# 3.78e-19
C2732 B15 a_4441_n1814# 0.2191f
C2733 B8 a_5288_n2068# 3.03e-19
C2734 A3 a_2273_n254# 0.037805f
C2735 a_798_n1194# a_143_n1036# 0.079554f
C2736 a_3832_n3674# a_2995_n4294# 1.4e-19
C2737 a_4000_n3674# a_3946_n2306# 7.6e-20
C2738 DVDD a_1557_46# 0.364955f
C2739 a_3946_n1066# a_3874_n2460# 0.002572f
C2740 a_3543_n342# a_5855_n574# 2.52e-19
C2741 a_3765_n600# a_4523_n574# 0.001897f
C2742 a_3669_n342# a_4691_n574# 2.26e-19
C2743 a_4204_n3054# a_4691_n2734# 5.41e-19
C2744 a_541_n3308# a_n131_n4294# 5.55e-19
C2745 a_3322_n4062# a_3904_n3674# 0.023518f
C2746 B1 a_1641_412# 0.020016f
C2747 A1 a_1997_412# 0.011819f
C2748 a_143_n2276# a_541_n3308# 6.58e-21
C2749 DVDD a_3736_412# 6.64e-19
C2750 Cin a_2254_46# 0.034155f
C2751 B6 a_101_n2434# 1.3e-19
C2752 DVDD a_2543_n254# 2.46e-19
C2753 a_636_n4294# a_n131_n3054# 0.003854f
C2754 a_5402_n2306# A8 0.780011f
C2755 A7 A11 0.006192f
C2756 a_3874_n1220# a_3322_n1582# 0.022847f
C2757 a_3736_n2068# a_3904_n2434# 0.007578f
C2758 a_3543_n342# a_3685_n1775# 9.8e-19
C2759 A7 a_1641_n2434# 1.4e-21
C2760 a_101_n2434# a_143_n3516# 0.008359f
C2761 B12 a_5402_174# 0.181244f
C2762 a_1557_46# a_1467_412# 0.006823f
C2763 A13 a_2908_n600# 2.15e-19
C2764 a_5402_n2306# a_5773_n1814# 5.92e-19
C2765 a_101_46# a_894_412# 4.35e-21
C2766 B1 a_n131_n1814# 2.07e-21
C2767 a_143_n2276# a_636_n1814# 0.030796f
C2768 a_636_n574# a_798_46# 0.012687f
C2769 a_3946_174# a_3322_n1582# 0.008526f
C2770 a_3874_20# a_6023_n574# 4.33e-19
C2771 a_143_n2276# B3 0.022193f
C2772 a_1261_n4320# a_1479_n3974# 0.007234f
C2773 a_3736_n2434# a_4000_n2434# 8.12e-20
C2774 a_4204_n574# a_4000_46# 7.87e-20
C2775 A1 a_1557_n1194# 2.88e-19
C2776 A7 a_2350_n3674# 5.43e-19
C2777 a_2995_n4294# a_4691_n1494# 4.48e-19
C2778 a_1557_n2434# a_3946_n2306# 0.001288f
C2779 a_5456_n3674# a_4204_n3054# 0.045338f
C2780 a_636_n3054# a_2995_n4294# 0.004323f
C2781 a_3322_n1582# a_4523_n574# 3.8e-19
C2782 a_798_n2434# a_894_n2434# 0.005587f
C2783 a_101_n3674# a_636_n4294# 0.201352f
C2784 a_5360_n2434# B10 1.22e-20
C2785 a_185_46# a_541_46# 0.008475f
C2786 a_2273_n2734# a_3322_n4062# 0.0099f
C2787 A13 a_3874_20# 0.512147f
C2788 B13 a_1557_46# 2.32e-20
C2789 a_3589_n1448# a_3434_n1546# 0.005193f
C2790 a_2254_n1194# a_2422_n828# 0.007578f
C2791 a_101_n1194# a_894_n1194# 3.78e-19
C2792 B13 a_3736_412# 3.18e-19
C2793 a_143_n2276# a_1291_n574# 7.74e-19
C2794 DVDD a_4000_412# 0.154852f
C2795 a_5192_46# a_5360_46# 0.00792f
C2796 A15 a_3765_n600# 1.85e-19
C2797 A6 a_541_n3674# 0.047225f
C2798 a_4000_n3674# a_4363_n3674# 0.008475f
C2799 a_2273_n254# a_1201_n574# 0.202439f
C2800 a_143_n1036# a_1201_n1814# 0.022242f
C2801 A3 a_1997_n828# 0.011819f
C2802 a_3874_n1220# a_3946_n1066# 0.287345f
C2803 a_101_n1194# a_143_n1036# 0.219575f
C2804 a_101_n2434# a_n131_n4294# 2.69e-19
C2805 a_1557_n2434# a_1201_n3054# 0.076462f
C2806 a_143_n2276# a_2783_n1775# 0.003083f
C2807 a_636_n3054# a_1201_n4294# 7.1e-20
C2808 a_5456_n3308# a_5402_n3546# 0.004108f
C2809 A1 a_1647_n574# 1.5e-19
C2810 a_3543_n2822# B10 0.057188f
C2811 a_143_n2276# a_101_n2434# 0.224993f
C2812 DVDD a_4363_n1194# 0.001386f
C2813 a_5402_n2306# a_4204_n3054# 0.008359f
C2814 B2 a_n131_n1814# 0.057188f
C2815 a_3434_n1546# a_3543_n2822# 1.28e-20
C2816 DVDD a_6153_n3308# 5.28e-19
C2817 B11 a_n131_n4294# 1.25e-20
C2818 Cin a_2350_n1194# 1.03e-20
C2819 DVDD A3 0.480085f
C2820 B11 a_143_n2276# 1.52e-20
C2821 a_3946_n1066# a_3946_174# 0.007318f
C2822 B9 a_3874_n3700# 1.11e-19
C2823 a_1201_n1814# a_2569_n1775# 1.29e-20
C2824 DVDD B9 0.594006f
C2825 a_5402_n1066# a_6153_n1194# 0.006958f
C2826 a_1557_n1194# a_2315_n1775# 0.027489f
C2827 a_636_n1814# a_1968_n1814# 1.72e-19
C2828 a_2422_n2068# a_n131_n1814# 4.28e-20
C2829 A15 a_3946_n2306# 2.88e-19
C2830 B8 a_5819_n1194# 8.1e-22
C2831 a_3736_n1194# a_2908_n600# 0.00792f
C2832 a_3874_20# a_5402_174# 0.172114f
C2833 a_4204_n574# a_5192_46# 1.96e-19
C2834 A2 a_1557_n1194# 0.001406f
C2835 B0 a_n41_n574# 0.056561f
C2836 a_3655_n1516# a_2273_n254# 2.2e-20
C2837 B3 a_1968_n1814# 0.002893f
C2838 a_5402_n2306# a_5360_n1194# 9.75e-22
C2839 DVDD a_3589_n3928# 2.55e-19
C2840 B4 a_185_n1194# 8.1e-22
C2841 a_3946_n2306# B8 3.07e-19
C2842 a_3874_n1220# a_4691_n574# 1.21e-19
C2843 a_2995_n4294# a_5288_n2068# 4.99e-19
C2844 B2 a_798_n1194# 0.078521f
C2845 a_3543_n342# a_6023_n2734# 2.42e-19
C2846 a_n131_n1814# a_315_n3054# 2.76e-19
C2847 a_3736_n2434# a_3904_n2434# 0.00792f
C2848 a_1557_n2434# a_636_n4294# 0.002601f
C2849 A10 a_5192_n3674# 7.66e-19
C2850 A15 a_3322_n1582# 0.037805f
C2851 A11 a_4691_n4294# 0.007493f
C2852 B13 a_4000_412# 0.005326f
C2853 A13 a_4363_412# 0.011562f
C2854 A6 a_1201_n4294# 1.6e-19
C2855 a_5402_n3546# a_5288_n3308# 4.35e-21
C2856 a_4204_n574# a_5456_n828# 0.087066f
C2857 a_4000_n1194# a_4363_n1194# 0.008475f
C2858 DVDD a_n41_n1814# 0.265726f
C2859 A2 a_147_n1494# 0.001052f
C2860 A11 a_3874_n3700# 0.51166f
C2861 a_3736_n2068# B9 3.18e-19
C2862 B1 a_1201_n1814# 6.28e-19
C2863 DVDD A11 0.470479f
C2864 a_5773_n1814# a_6023_n574# 3.47e-20
C2865 a_5456_n3308# a_5288_n3308# 2.18e-19
C2866 a_3946_174# a_2254_46# 2.97e-20
C2867 A9 a_4000_n2434# 0.046632f
C2868 DVDD a_1641_n2434# 0.001386f
C2869 a_3874_n2460# A5 2.02e-20
C2870 B13 a_4363_n1194# 2.95e-21
C2871 a_3765_n3080# a_2543_n2734# 1.71e-20
C2872 a_3669_n2822# a_3627_n2734# 0.008516f
C2873 a_636_n574# a_1997_412# 0.112124f
C2874 a_3434_n4026# a_4441_n4294# 0.053796f
C2875 a_3434_n4026# a_3861_n3080# 5.85e-21
C2876 a_4441_n4294# a_3669_n2822# 0.188936f
C2877 a_636_n3054# a_2315_n1775# 8.78e-19
C2878 a_5773_n4294# a_3543_n2822# 0.188784f
C2879 a_1557_n2434# a_1261_n1840# 1.81e-19
C2880 a_3655_n3996# a_3765_n3080# 2.4e-19
C2881 B2 a_315_n1814# 0.007771f
C2882 A2 B4 1.32e-19
C2883 a_3669_n2822# a_3861_n3080# 0.006573f
C2884 DVDD a_4523_n3054# 0.005567f
C2885 a_n131_n574# a_2254_n1194# 3.29e-19
C2886 a_1201_n1814# a_1641_n828# 3.93e-19
C2887 B15 a_3543_n342# 0.00432f
C2888 a_2254_n3674# a_n131_n3054# 3.29e-19
C2889 a_636_n1814# a_1467_n828# 7.45e-20
C2890 a_3765_n600# a_3861_n600# 0.197466f
C2891 DVDD a_1201_n574# 0.179937f
C2892 a_n71_n600# a_1201_n574# 2.84e-19
C2893 A5 a_n131_n3054# 0.022989f
C2894 B3 a_1467_n828# 4.23e-20
C2895 a_3669_n2822# a_3904_n2434# 3.97e-19
C2896 B2 A4 1.23e-19
C2897 a_n41_n3054# a_n71_n3080# 0.025037f
C2898 B10 a_5855_n4294# 0.007771f
C2899 a_3946_n1066# A15 0.791917f
C2900 B15 a_4441_n574# 7.54e-19
C2901 a_5402_n1066# a_5456_n828# 0.004108f
C2902 a_3946_n3546# B10 3.07e-19
C2903 a_1997_46# a_2254_46# 0.023012f
C2904 a_3368_n3928# a_3226_n4062# 0.007833f
C2905 a_2497_n4255# a_1968_n4294# 4.9e-19
C2906 B12 a_5456_46# 0.005557f
C2907 A12 a_5819_46# 0.050725f
C2908 a_4441_n4294# A9 8.18e-21
C2909 a_185_n828# a_n131_n1814# 5.74e-19
C2910 B2 a_1201_n1814# 4.1e-19
C2911 a_2995_n4294# a_3765_n600# 5.32e-19
C2912 B2 a_101_n1194# 0.181244f
C2913 A9 a_3861_n3080# 0.022989f
C2914 B14 a_5192_n828# 3.18e-19
C2915 a_1557_46# a_3904_46# 2.97e-20
C2916 a_1997_n3308# a_636_n4294# 0.112124f
C2917 a_3874_20# a_3832_412# 1.35e-20
C2918 a_541_n2068# a_894_n2068# 2.18e-19
C2919 DVDD a_3655_n1516# 0.194591f
C2920 a_1261_n4320# a_1261_n3080# 0.002078f
C2921 a_n71_n4320# a_n131_n3054# 1.01e-20
C2922 a_5360_n3674# B10 0.078521f
C2923 a_3904_46# a_3736_412# 0.007578f
C2924 a_4000_n828# a_2908_n600# 0.023311f
C2925 a_3736_n828# a_3669_n342# 1.98e-19
C2926 Cin a_n131_n4294# 0.001045f
C2927 a_2254_n2434# a_1557_n1194# 1.25e-21
C2928 Cin a_143_n2276# 0.02168f
C2929 A15 a_4691_n574# 7.81e-20
C2930 B6 a_n131_n3054# 7.86e-19
C2931 a_3322_n1582# a_3861_n600# 0.158736f
C2932 A9 a_3904_n2434# 0.114466f
C2933 a_6023_n254# a_3543_n342# 6.93e-20
C2934 a_4204_n574# a_3765_n600# 0.068052f
C2935 a_2995_n4294# a_5819_n1194# 1.55e-21
C2936 a_5819_n2068# B14 5.74e-19
C2937 a_636_n574# a_1647_n574# 2.35e-19
C2938 a_3832_n3674# a_3904_n3674# 0.005587f
C2939 DVDD a_5855_n1814# 0.008551f
C2940 a_3177_n1814# a_3543_n342# 0.002372f
C2941 a_1479_n2734# a_1201_n3054# 0.004527f
C2942 a_143_n3516# a_n131_n3054# 0.182595f
C2943 a_2273_n2734# a_1261_n3080# 6.57e-19
C2944 a_143_n1036# a_798_46# 0.0021f
C2945 a_3946_n2306# a_2995_n4294# 0.113366f
C2946 a_3874_n2460# a_5402_n2306# 0.172114f
C2947 B9 a_3736_n2434# 6.11e-20
C2948 a_5402_n2306# a_6153_n2434# 0.006958f
C2949 a_3322_n4062# a_4523_n4294# 3.9e-20
C2950 a_4204_n574# a_5819_n1194# 0.033252f
C2951 B6 a_894_n3308# 2.91e-19
C2952 a_1557_46# a_2363_n254# 6.28e-19
C2953 a_n71_n4320# a_101_n3674# 0.003994f
C2954 a_5773_n4294# a_5855_n4294# 0.006406f
C2955 a_2995_n4294# a_3322_n1582# 0.014561f
C2956 a_5192_n3308# B10 3.18e-19
C2957 B6 a_101_n3674# 0.181244f
C2958 a_143_n3516# a_894_n3308# 2.9e-19
C2959 a_1557_n3674# a_3322_n4062# 8.35e-21
C2960 a_2273_n2734# a_798_n3674# 2.74e-19
C2961 B7 a_1647_n4294# 0.007771f
C2962 a_2995_n4294# a_1201_n3054# 0.004827f
C2963 a_4441_n4294# a_5402_n3546# 0.005934f
C2964 a_966_n3674# a_798_n3674# 0.00792f
C2965 a_143_n2276# a_3874_n2460# 1.28e-20
C2966 a_3861_n3080# a_5402_n3546# 2.05e-19
C2967 a_1997_n2068# a_1557_n2434# 0.004411f
C2968 a_4441_n3054# a_3946_n3546# 1.81e-19
C2969 a_101_n3674# a_143_n3516# 0.219575f
C2970 A0 a_1261_n600# 6.77e-21
C2971 a_2254_n2434# a_636_n3054# 0.062548f
C2972 B0 a_n71_n600# 0.226175f
C2973 DVDD B0 0.775788f
C2974 a_3904_46# a_4000_412# 0.02283f
C2975 B5 a_n71_n3080# 3.52e-21
C2976 a_3322_n1582# a_4204_n574# 0.01799f
C2977 a_2254_n3674# a_1557_n2434# 4.59e-21
C2978 DVDD a_147_n3974# 0.001263f
C2979 a_5360_n2434# a_5288_n2434# 0.005587f
C2980 DVDD a_5773_n3054# 0.172232f
C2981 a_894_n3674# a_101_n3674# 3.78e-19
C2982 S15 a_143_n2276# 9.71e-19
C2983 a_1291_n1814# B5 2.83e-19
C2984 a_1557_n1194# B15 2.32e-20
C2985 a_1557_n2434# A5 0.792469f
C2986 a_3946_n1066# a_3861_n600# 6.4e-19
C2987 a_2273_n254# a_2908_n600# 2.31e-19
C2988 a_1997_n2434# a_2422_n2434# 8.12e-20
C2989 A3 a_1641_n1194# 0.051667f
C2990 a_1997_n3674# a_2350_n3674# 2.18e-19
C2991 a_798_n1194# a_1467_n1194# 5.49e-20
C2992 Cin a_1968_n1814# 0.299183f
C2993 a_n131_n3054# a_n131_n4294# 0.001745f
C2994 a_1201_n3054# a_1201_n4294# 0.15552f
C2995 B11 a_4000_n3308# 0.005326f
C2996 a_185_412# a_541_412# 0.009846f
C2997 a_143_n2276# a_n131_n3054# 0.003969f
C2998 DVDD a_4363_n2068# 0.160791f
C2999 B1 a_798_46# 2.55e-19
C3000 Cin a_966_412# 2.78e-19
C3001 a_185_n2068# a_n131_n1814# 0.003904f
C3002 B9 a_3669_n2822# 6.28e-19
C3003 a_5402_174# a_5360_n1194# 1.16e-19
C3004 a_1467_n2068# DVDD 4.94e-19
C3005 a_2995_n4294# a_636_n4294# 0.004633f
C3006 a_3543_n342# a_2569_n1775# 7.26e-19
C3007 a_5402_174# a_5288_412# 4.35e-21
C3008 a_3589_n3928# a_3434_n4026# 0.005193f
C3009 a_3736_n3308# a_3322_n4062# 1.91e-19
C3010 a_5402_n1066# a_5819_n1194# 0.067562f
C3011 a_3589_n3928# a_3669_n2822# 6.39e-19
C3012 a_894_n828# a_2273_n254# 1.6e-20
C3013 a_4363_n3674# a_2995_n4294# 8.14e-19
C3014 a_3946_n1066# a_2995_n4294# 0.008944f
C3015 a_3874_n1220# a_5402_n2306# 8.25e-20
C3016 a_185_n828# a_101_n1194# 0.030161f
C3017 a_1261_n4320# a_636_n3054# 9.91e-21
C3018 a_3861_n600# a_4691_n574# 0.058037f
C3019 a_894_n3308# a_n131_n4294# 3.32e-20
C3020 a_4204_n3054# a_4000_n3308# 5.14e-19
C3021 a_3322_n4062# a_4363_n3308# 0.001272f
C3022 DVDD a_3711_n254# 1.88e-19
C3023 Cin A13 1.35e-19
C3024 A9 a_4363_n1194# 1.4e-21
C3025 DVDD B12 0.746279f
C3026 a_636_n4294# a_1201_n4294# 0.105485f
C3027 a_101_n3674# a_n131_n4294# 0.034089f
C3028 B3 B5 0.004788f
C3029 B15 a_4691_n1494# 0.002951f
C3030 a_3832_n2068# a_4000_n2068# 2.18e-19
C3031 a_3946_n1066# a_4204_n574# 0.005791f
C3032 a_3669_n342# a_4523_n1814# 0.002223f
C3033 a_5402_n1066# a_3322_n1582# 5.68e-21
C3034 a_5773_n574# a_6023_n574# 0.025037f
C3035 A11 a_3434_n4026# 0.00356f
C3036 a_1557_n2434# a_143_n3516# 0.057421f
C3037 a_636_n3054# a_2273_n2734# 3.49e-19
C3038 A11 a_3669_n2822# 0.077871f
C3039 A9 B9 1.25311f
C3040 A13 a_3669_n342# 0.001673f
C3041 a_1968_n4294# a_3322_n4062# 1.42e-19
C3042 a_2995_n4294# a_4691_n574# 4.81e-19
C3043 a_1291_n1814# a_2273_n254# 1.57e-19
C3044 a_143_n1036# a_1997_412# 1.25e-20
C3045 B2 a_798_46# 1.22e-20
C3046 a_3322_n1582# a_2315_n1775# 2.2e-20
C3047 a_636_n4294# a_1467_n3308# 7.45e-20
C3048 a_1968_n4294# a_1479_n3974# 3.05e-19
C3049 A6 a_1261_n4320# 6.77e-21
C3050 a_1997_n1194# a_2350_n1194# 2.18e-19
C3051 a_1997_n3308# a_2254_n3674# 0.02283f
C3052 a_4523_n3054# a_3669_n2822# 1.02e-20
C3053 A13 a_5773_n574# 1.38e-21
C3054 a_1997_n1194# A5 6.84e-21
C3055 a_1997_n3308# A5 8.69e-21
C3056 a_n131_n3054# a_1968_n1814# 4.03e-21
C3057 a_1201_n3054# a_2315_n1775# 2.07e-19
C3058 a_798_n2434# a_1467_n2434# 5.49e-20
C3059 a_143_n2276# a_n71_n1840# 7.64e-19
C3060 a_2995_n4294# a_3368_n1775# 6.81e-19
C3061 a_1647_n1814# a_1261_n1840# 0.006406f
C3062 A0 a_541_46# 0.047225f
C3063 B0 a_185_46# 0.021045f
C3064 DVDD a_894_46# 8.89e-20
C3065 a_4204_n574# a_4691_n574# 0.016475f
C3066 a_2908_n600# a_1997_n828# 9.34e-20
C3067 a_n131_n1814# a_2254_n1194# 0.008425f
C3068 a_1467_n1194# a_1201_n1814# 9.84e-21
C3069 a_101_n2434# B5 7.19e-19
C3070 a_636_n1814# a_966_n1194# 3.15e-19
C3071 DVDD a_2908_n600# 0.834969f
C3072 A6 a_2273_n2734# 5.21e-20
C3073 A11 A9 0.002462f
C3074 A4 a_185_n2068# 0.011602f
C3075 a_3322_n1582# a_3685_n1775# 0.005265f
C3076 A1 a_1261_n1840# 8.18e-21
C3077 A6 a_966_n3674# 7.66e-19
C3078 B13 B12 0.003904f
C3079 a_101_46# a_541_n1194# 4.36e-20
C3080 a_3946_n1066# a_5402_n1066# 0.003292f
C3081 a_1557_n2434# a_n131_n4294# 7.63e-19
C3082 a_636_n1814# a_2273_n254# 0.022847f
C3083 a_6153_n3308# a_5402_n3546# 0.006823f
C3084 a_1557_n1194# a_143_n1036# 0.005791f
C3085 a_143_n2276# a_1557_n2434# 0.095682f
C3086 A9 a_4523_n3054# 1.5e-19
C3087 A14 a_4441_n1814# 6.77e-21
C3088 a_3655_n1516# a_3669_n2822# 3.16e-19
C3089 DVDD a_894_n828# 5.34e-19
C3090 B3 a_2273_n254# 0.040998f
C3091 a_5402_174# a_5773_n574# 0.003994f
C3092 DVDD a_3874_20# 0.895778f
C3093 a_1557_46# a_1261_n600# 0.002379f
C3094 A0 a_1557_46# 0.001406f
C3095 a_3655_n1516# a_3904_46# 7.07e-21
C3096 a_5402_174# a_5456_n1194# 4.36e-20
C3097 Cin a_2350_412# 2.58e-19
C3098 B1 a_1997_412# 0.005326f
C3099 A1 a_2254_46# 0.114466f
C3100 a_1557_n1194# a_2569_n1775# 4.55e-19
C3101 a_3736_n1194# a_3669_n342# 5.8e-19
C3102 a_4000_n1194# a_2908_n600# 0.023012f
C3103 DVDD a_5456_n2434# 8.16e-19
C3104 a_1997_n3308# a_143_n3516# 5.14e-19
C3105 a_2363_n254# a_1201_n574# 0.006083f
C3106 DVDD a_2783_n4255# 0.001765f
C3107 B7 A11 2.72e-20
C3108 A7 B11 2.72e-20
C3109 a_5402_n2306# B8 0.181244f
C3110 A15 a_3736_n828# 1.05e-19
C3111 a_6023_n1814# A14 0.007489f
C3112 B7 a_1641_n2434# 3.27e-20
C3113 A5 a_1479_n2734# 9.63e-19
C3114 a_143_n1036# a_1647_n574# 0.003613f
C3115 a_2273_n254# a_1291_n574# 5.44e-19
C3116 a_1557_n3674# a_1261_n3080# 1.81e-19
C3117 a_4000_n2434# a_3904_n2434# 0.023012f
C3118 A10 a_5456_n3674# 0.047225f
C3119 B13 a_2908_n600# 6.76e-20
C3120 a_n71_n1840# a_1968_n1814# 1.26e-20
C3121 DVDD a_n71_n3080# 0.177213f
C3122 A2 a_1261_n1840# 6.77e-21
C3123 a_4204_n574# a_6153_n828# 1.23e-20
C3124 A9 a_3655_n1516# 0.002599f
C3125 DVDD a_1291_n1814# 0.259614f
C3126 a_2273_n254# a_2783_n1775# 0.006879f
C3127 a_143_n2276# A15 1.11e-19
C3128 a_1997_n2068# a_2995_n4294# 5.63e-19
C3129 a_2254_n2434# a_3946_n2306# 2.97e-20
C3130 A11 a_5402_n3546# 1.36e-19
C3131 a_2254_n3674# a_2995_n4294# 0.005991f
C3132 A13 a_3874_n1220# 0.004204f
C3133 a_1557_n3674# a_798_n3674# 0.031298f
C3134 B1 a_1557_n1194# 3.5e-19
C3135 B7 a_2350_n3674# 7.33e-20
C3136 a_2995_n4294# A5 0.00648f
C3137 a_3669_n2822# a_3795_n2734# 1.46e-22
C3138 a_3765_n3080# a_3711_n2734# 0.009339f
C3139 a_3543_n2822# a_3322_n4062# 0.034265f
C3140 a_3946_n2306# a_3904_n3674# 4.59e-21
C3141 a_2995_n4294# a_4691_n2734# 4.8e-19
C3142 DVDD a_541_n3308# 0.157566f
C3143 B13 a_3874_20# 1.25937f
C3144 a_2254_46# a_2315_n1775# 7.07e-21
C3145 A13 a_3946_174# 0.792469f
C3146 a_4441_n4294# a_3861_n3080# 9.27e-21
C3147 a_1557_n2434# a_1968_n1814# 5.1e-20
C3148 A10 a_5402_n2306# 0.003407f
C3149 DVDD a_4363_412# 0.160791f
C3150 a_3765_n3080# a_4441_n3054# 0.243071f
C3151 a_5288_46# a_5360_46# 0.005587f
C3152 DVDD a_5855_n3054# 0.005567f
C3153 a_2254_n2434# a_1201_n3054# 4.74e-19
C3154 a_5288_n3674# a_5456_n3674# 2.18e-19
C3155 a_1201_n1814# a_2254_n1194# 0.023649f
C3156 B15 a_3765_n600# 0.00216f
C3157 B6 a_541_n3674# 0.005557f
C3158 a_2254_n3674# a_1201_n4294# 0.023649f
C3159 a_636_n1814# a_1997_n828# 0.112124f
C3160 a_1557_n1194# a_1641_n828# 0.030161f
C3161 a_1997_n1194# a_143_n2276# 0.001591f
C3162 a_1997_n3308# a_143_n2276# 5.5e-19
C3163 a_3322_n1582# a_3904_n3674# 5.66e-21
C3164 a_1479_n2734# a_143_n3516# 5.41e-19
C3165 A13 a_4523_n574# 1.5e-19
C3166 B3 a_1997_n828# 0.005326f
C3167 a_3861_n3080# a_3904_n2434# 3.5e-19
C3168 A5 a_1201_n4294# 0.001673f
C3169 B1 a_1647_n574# 0.007771f
C3170 DVDD a_636_n1814# 1.04236f
C3171 a_n41_n3054# a_n131_n3054# 0.131556f
C3172 a_541_n3674# a_143_n3516# 0.045338f
C3173 B14 a_3434_n1546# 1.57e-20
C3174 DVDD B3 0.619467f
C3175 a_541_n3674# a_894_n3674# 2.18e-19
C3176 A3 a_1261_n600# 1.75e-19
C3177 a_5402_n1066# a_6153_n828# 0.006823f
C3178 a_1997_n3308# a_1641_n3308# 0.009846f
C3179 a_2783_n4255# a_2569_n4255# 0.005572f
C3180 DVDD A8 0.480037f
C3181 B15 a_3946_n2306# 3.5e-19
C3182 a_3946_174# a_5402_174# 0.003292f
C3183 A9 a_5773_n3054# 1.38e-21
C3184 B2 a_1557_n1194# 3.07e-19
C3185 a_2995_n4294# a_143_n3516# 0.001341f
C3186 a_4204_n574# a_5288_46# 1.66e-19
C3187 a_2350_n3308# a_636_n4294# 1.35e-20
C3188 DVDD a_5773_n1814# 0.190735f
C3189 Cin a_n41_n574# 1.35e-19
C3190 a_798_n2434# a_966_n2068# 0.007578f
C3191 B0 a_315_n574# 0.007771f
C3192 a_1261_n4320# a_1201_n3054# 7.34e-21
C3193 a_n71_n4320# a_1201_n4294# 3.93e-19
C3194 a_2315_n4255# a_n131_n3054# 5.6e-20
C3195 a_5819_n3308# B10 0.033026f
C3196 DVDD a_1291_n574# 0.238543f
C3197 a_4000_n828# a_3669_n342# 4.28e-19
C3198 a_636_n574# a_1261_n1840# 9.91e-21
C3199 a_636_n4294# a_3904_n3674# 2.15e-20
C3200 Cin a_3368_n1448# 3.11e-19
C3201 B15 a_3322_n1582# 0.040998f
C3202 B11 a_4691_n4294# 0.056553f
C3203 B6 a_1201_n4294# 4.1e-19
C3204 B13 a_4363_412# 0.020016f
C3205 a_894_n2434# A4 5.43e-19
C3206 a_6023_n254# a_3765_n600# 2.05e-20
C3207 A9 a_4363_n2068# 0.011562f
C3208 a_4691_n254# a_3861_n600# 9.28e-20
C3209 a_1479_n1494# a_1201_n1814# 0.002666f
C3210 DVDD a_2783_n1775# 0.001765f
C3211 DVDD a_101_n2434# 0.394947f
C3212 B11 a_3874_n3700# 1.25417f
C3213 B2 a_147_n1494# 0.002402f
C3214 a_143_n3516# a_1201_n4294# 0.022242f
C3215 a_2273_n2734# a_1201_n3054# 0.202439f
C3216 a_3589_n1448# a_3543_n342# 0.001075f
C3217 a_5360_n2434# a_3543_n342# 0.00219f
C3218 a_2995_n4294# a_5402_n2306# 0.224913f
C3219 a_143_n2276# a_1479_n2734# 2.75e-19
C3220 a_541_n3674# a_n131_n4294# 0.001186f
C3221 DVDD B11 0.610099f
C3222 B9 a_4000_n2434# 0.005557f
C3223 a_3874_n2460# B5 2.79e-20
C3224 a_2995_n4294# a_3736_n828# 3.11e-20
C3225 a_636_n574# a_2254_46# 0.062548f
C3226 a_4204_n3054# a_4691_n4294# 1.59e-20
C3227 A13 A15 0.002462f
C3228 a_1557_46# a_2543_n254# 3.01e-19
C3229 a_1261_n4320# a_636_n4294# 0.015611f
C3230 A5 a_2315_n1775# 0.002599f
C3231 B2 B4 0.008756f
C3232 a_2273_n2734# a_966_n3308# 1.79e-20
C3233 a_3946_n3546# a_3322_n4062# 0.142863f
C3234 a_143_n3516# a_1467_n3308# 5.15e-20
C3235 a_3874_n3700# a_4204_n3054# 0.026336f
C3236 a_2790_n1448# a_3434_n1546# 8.12e-20
C3237 a_3543_n2822# a_3543_n342# 3.71e-20
C3238 a_3322_n1582# a_3832_n828# 2.27e-19
C3239 A14 a_3543_n342# 0.02685f
C3240 a_2995_n4294# a_n131_n4294# 0.022241f
C3241 a_143_n2276# a_2995_n4294# 0.202092f
C3242 A6 a_1557_n3674# 0.001406f
C3243 DVDD a_4204_n3054# 0.780566f
C3244 a_636_n4294# a_2273_n2734# 0.022847f
C3245 a_2350_n2068# a_1557_n2434# 4.35e-21
C3246 Cin a_2273_n254# 0.056021f
C3247 a_5773_n3054# a_5402_n3546# 5.92e-19
C3248 a_1261_n600# a_1201_n574# 0.243071f
C3249 A0 a_1201_n574# 4.94e-20
C3250 B5 a_n131_n3054# 0.033034f
C3251 a_4204_n574# a_4691_n254# 5.41e-19
C3252 a_5360_n3674# a_3322_n4062# 2.74e-19
C3253 a_966_n3674# a_636_n4294# 3.15e-19
C3254 a_3946_n1066# B15 0.175017f
C3255 B11 a_3832_n3308# 2.91e-19
C3256 B4 a_315_n3054# 0.007771f
C3257 A11 a_4000_n2434# 6.84e-21
C3258 a_2273_n254# a_3669_n342# 6.64e-20
C3259 a_3177_n1814# a_3322_n1582# 0.00841f
C3260 a_636_n3054# a_315_n3054# 3.68e-19
C3261 a_798_n2434# a_n131_n1814# 0.00219f
C3262 A14 a_5288_n1194# 5.43e-19
C3263 DVDD a_5360_n1194# 0.234243f
C3264 a_2995_n4294# a_1641_n3308# 5.59e-19
C3265 a_2350_46# a_2254_46# 0.005587f
C3266 B12 a_5819_46# 0.021045f
C3267 B11 a_4697_n3308# 4.23e-20
C3268 a_1201_n4294# a_n131_n4294# 1.11131f
C3269 a_143_n2276# a_1201_n4294# 0.01677f
C3270 a_4441_n4294# B9 3.66e-21
C3271 DVDD a_5192_n2068# 6.64e-19
C3272 DVDD a_5288_412# 5.1e-19
C3273 a_541_n828# a_n131_n1814# 5.55e-19
C3274 a_1647_n1814# a_143_n2276# 0.002427f
C3275 a_541_n2434# a_101_n2434# 0.044963f
C3276 B9 a_3861_n3080# 0.033034f
C3277 a_3946_174# a_3832_412# 4.35e-21
C3278 a_3874_20# a_3904_46# 0.062548f
C3279 A14 a_5819_n2434# 1.15e-19
C3280 a_4000_412# a_3736_412# 1.31e-19
C3281 a_3832_n2068# a_3322_n4062# 1.21e-20
C3282 a_3832_n3308# a_4204_n3054# 1.19e-20
C3283 A1 a_143_n2276# 0.001332f
C3284 A7 a_n131_n3054# 3.72e-19
C3285 B9 a_3904_n2434# 0.077428f
C3286 a_5402_n1066# a_5402_n2306# 0.002006f
C3287 B15 a_4691_n574# 0.001447f
C3288 a_3861_n600# a_6023_n574# 0.131556f
C3289 a_1641_n3308# a_1201_n4294# 3.93e-19
C3290 a_4204_n3054# a_4697_n3308# 5.15e-20
C3291 a_3322_n4062# a_5192_n3308# 1.79e-20
C3292 a_143_n2276# a_1467_n3308# 6.47e-21
C3293 a_541_n828# a_798_n1194# 0.02283f
C3294 a_3736_n1194# A15 7.66e-19
C3295 a_3946_n1066# a_3832_n828# 4.35e-21
C3296 a_3874_n1220# a_4000_n828# 0.112124f
C3297 A3 a_1557_46# 3.41e-19
C3298 a_143_n2276# a_185_n1194# 1.55e-21
C3299 S15 a_2273_n254# 0.002239f
C3300 a_143_n1036# a_894_412# 3.3e-20
C3301 a_3946_174# a_4000_n828# 5.56e-19
C3302 A11 a_4441_n4294# 0.084607f
C3303 a_1557_n2434# a_2363_n2734# 6.28e-19
C3304 A11 a_3861_n3080# 3.72e-19
C3305 A13 a_3861_n600# 0.022989f
C3306 a_3226_n4062# a_3322_n4062# 0.318695f
C3307 A13 a_5360_46# 0.001236f
C3308 A7 a_101_n3674# 1.36e-19
C3309 a_1997_n2068# a_2254_n2434# 0.02283f
C3310 a_n41_n574# a_n71_n1840# 3.47e-20
C3311 a_3322_n1582# a_2569_n1775# 3.13e-19
C3312 Cin a_1997_n828# 1.3e-19
C3313 a_185_n1194# a_541_n1194# 0.008475f
C3314 a_1997_n3308# a_2422_n3308# 1.31e-19
C3315 a_2254_n3674# a_2350_n3308# 0.004869f
C3316 A11 a_3904_n2434# 1.29e-20
C3317 a_4523_n3054# a_3861_n3080# 0.005159f
C3318 a_4691_n3054# a_3765_n3080# 0.074717f
C3319 a_6023_n3054# a_3543_n2822# 4.81e-19
C3320 a_5456_n2068# A8 0.011819f
C3321 a_2254_n2434# A5 0.114466f
C3322 a_1201_n4294# a_1968_n1814# 3.6e-19
C3323 DVDD Cin 1.08579f
C3324 A0 B0 1.27934f
C3325 A1 a_1479_n254# 9.63e-19
C3326 Cin a_n71_n600# 1.52e-19
C3327 a_2995_n4294# a_4523_n1814# 0.001631f
C3328 a_143_n2276# a_2315_n1775# 0.011235f
C3329 a_2254_n3674# a_3904_n3674# 0.004465f
C3330 a_4204_n574# a_6023_n574# 0.002038f
C3331 a_3543_n342# a_2254_n1194# 1.02e-19
C3332 a_2908_n600# a_2350_n828# 2.04e-20
C3333 a_11_n3308# a_n131_n1814# 4.61e-21
C3334 a_1557_n2434# a_2350_n2434# 3.53e-19
C3335 A2 a_143_n2276# 2.96e-19
C3336 a_798_n2434# A4 0.114467f
C3337 a_3736_n3674# a_3669_n2822# 5.8e-19
C3338 A13 a_2995_n4294# 3.87e-19
C3339 a_1557_n1194# a_1467_n1194# 0.006958f
C3340 a_636_n1814# a_1641_n1194# 0.033252f
C3341 a_1557_n2434# B5 0.17279f
C3342 DVDD a_3669_n342# 0.365382f
C3343 B3 a_1641_n1194# 0.019568f
C3344 a_5402_174# a_3861_n600# 0.004436f
C3345 Cin a_1467_412# 4.69e-20
C3346 a_2995_n4294# a_3685_n4255# 6.59e-20
C3347 A13 a_4204_n574# 0.051784f
C3348 a_5773_n4294# B10 0.226175f
C3349 A14 a_6153_n1194# 4.78e-19
C3350 a_3874_n1220# a_2273_n254# 1.14e-21
C3351 a_143_n2276# a_3685_n1775# 2.28e-19
C3352 a_5402_174# a_5360_46# 0.057724f
C3353 a_798_n2434# a_101_n1194# 1.25e-21
C3354 DVDD a_5773_n574# 0.171897f
C3355 A2 a_541_n1194# 0.047225f
C3356 DVDD a_5456_n1194# 8.16e-19
C3357 a_3655_n1516# a_3861_n3080# 6e-20
C3358 a_4441_n1814# a_3765_n3080# 5.51e-20
C3359 a_3874_n2460# a_3874_n3700# 8.69e-20
C3360 a_966_n828# a_2273_n254# 1.79e-20
C3361 a_3322_n4062# a_3832_n2434# 6.08e-20
C3362 a_1261_n4320# A5 8.18e-21
C3363 a_541_n828# a_101_n1194# 0.004108f
C3364 a_1557_46# a_1201_n574# 0.076462f
C3365 DVDD a_3874_n2460# 0.912323f
C3366 a_5402_n3546# a_5456_n2434# 1.67e-20
C3367 a_3832_n2068# a_3543_n342# 2.73e-20
C3368 a_143_n1036# a_1261_n1840# 5.74e-19
C3369 A7 a_1557_n2434# 3.41e-19
C3370 a_n131_n4294# a_3368_n4255# 3.93e-20
C3371 a_3655_n1516# a_3904_n2434# 4e-19
C3372 a_4000_n1194# a_3669_n342# 0.001261f
C3373 a_2254_n3674# a_2273_n2734# 0.023518f
C3374 a_2350_n3308# a_143_n3516# 1.19e-20
C3375 DVDD a_6153_n2434# 2.33e-19
C3376 a_2543_n254# a_1201_n574# 3.31e-19
C3377 a_2459_n254# a_1201_n1814# 0.001239f
C3378 DVDD S15 0.178784f
C3379 B9 a_4363_n1194# 3.27e-20
C3380 A1 A13 0.006192f
C3381 Cin B13 1.52e-20
C3382 DVDD a_6023_n3974# 5.73e-19
C3383 a_4691_n1814# a_4441_n3054# 9.75e-20
C3384 A15 a_4000_n828# 0.011819f
C3385 B11 a_3434_n4026# 0.002893f
C3386 A5 a_2273_n2734# 4.12e-19
C3387 a_1557_n3674# a_1201_n3054# 5.07e-20
C3388 A10 a_6153_n3674# 4.78e-19
C3389 A9 A8 0.019542f
C3390 B11 a_3669_n2822# 0.081283f
C3391 B13 a_3669_n342# 6.28e-19
C3392 a_2315_n1775# a_1968_n1814# 0.153192f
C3393 DVDD a_n131_n3054# 1.68115f
C3394 a_5402_174# a_4204_n574# 0.008359f
C3395 a_2350_n2068# a_2995_n4294# 5.05e-20
C3396 a_541_n2068# a_101_n2434# 0.004108f
C3397 a_3736_n1194# a_2995_n4294# 1.21e-19
C3398 a_2422_n3308# a_2995_n4294# 7.14e-20
C3399 B13 a_5773_n574# 3.52e-21
C3400 a_3655_n3996# a_3322_n4062# 0.236061f
C3401 a_3434_n4026# a_4204_n3054# 8.25e-20
C3402 a_143_n2276# a_636_n574# 2.79e-19
C3403 a_185_n2068# B4 0.033026f
C3404 a_5456_n2068# a_5192_n2068# 1.31e-19
C3405 a_5360_n2434# a_5288_n2068# 0.004869f
C3406 A0 a_894_46# 5.43e-19
C3407 Cin a_185_46# 0.033252f
C3408 DVDD a_966_46# 9.02e-20
C3409 a_3765_n3080# a_3322_n4062# 0.202439f
C3410 a_3669_n2822# a_4204_n3054# 0.022242f
C3411 B0 a_541_46# 0.005557f
C3412 a_1261_n4320# a_143_n3516# 5.74e-19
C3413 a_2995_n4294# a_4000_n3308# 0.001596f
C3414 DVDD a_894_n3308# 5.34e-19
C3415 a_3832_n1194# a_3322_n1582# 4.97e-19
C3416 a_636_n4294# a_1557_n3674# 0.287345f
C3417 B6 a_2273_n2734# 2.25e-20
C3418 a_n131_n574# a_n131_n1814# 0.001745f
C3419 a_1261_n600# a_2908_n600# 4.29e-21
C3420 a_3861_n3080# a_5773_n3054# 0.211818f
C3421 DVDD a_101_n3674# 0.391065f
C3422 a_5456_n3674# a_5819_n3674# 0.008475f
C3423 B1 a_1261_n1840# 3.66e-21
C3424 a_1201_n1814# a_2422_n828# 1.98e-19
C3425 A11 B9 0.007762f
C3426 B11 A9 0.004004f
C3427 B6 a_966_n3674# 6.11e-20
C3428 a_2254_n2434# a_143_n2276# 0.041493f
C3429 A12 B12 1.27934f
C3430 a_2422_n3308# a_1201_n4294# 1.98e-19
C3431 a_2422_n1194# a_143_n2276# 1.87e-19
C3432 a_1557_n1194# a_2254_n1194# 0.051953f
C3433 a_636_n1814# a_2350_n828# 1.35e-20
C3434 A6 a_n41_n4294# 0.007489f
C3435 a_4000_n3674# a_3874_n3700# 0.045338f
C3436 a_3832_n3674# a_3946_n3546# 2.79e-19
C3437 a_2350_n3308# a_143_n2276# 2.39e-20
C3438 A14 a_5456_n828# 0.011819f
C3439 a_143_n3516# a_2273_n2734# 0.01799f
C3440 B3 a_2350_n828# 2.91e-19
C3441 DVDD a_4000_n3674# 8.16e-19
C3442 DVDD a_3874_n1220# 1.03962f
C3443 a_1291_n3054# a_n131_n3054# 0.058037f
C3444 a_1647_n3054# a_1261_n3080# 0.006406f
C3445 a_966_n3674# a_143_n3516# 1.32e-19
C3446 a_n131_n4294# a_3904_n3674# 1.02e-19
C3447 a_2315_n4255# a_2995_n4294# 0.003116f
C3448 a_143_n2276# a_3904_n3674# 1.26e-19
C3449 B9 a_4523_n3054# 0.007771f
C3450 DVDD a_966_n828# 7.01e-19
C3451 A3 a_1201_n574# 1.85e-19
C3452 A8 a_5402_n3546# 6.66e-20
C3453 a_5402_n1066# a_5402_174# 0.007891f
C3454 A7 a_1997_n3308# 0.011819f
C3455 DVDD a_3946_174# 0.36446f
C3456 B0 a_1557_46# 3.07e-19
C3457 a_3434_n1546# a_n131_n1814# 2.79e-19
C3458 A9 a_4204_n3054# 0.051784f
C3459 a_3226_n1582# a_2908_n600# 1.21e-19
C3460 B1 a_2254_46# 0.077428f
C3461 Cin a_2422_412# 2.6e-19
C3462 DVDD a_101_46# 0.392196f
C3463 a_101_46# a_n71_n600# 0.003994f
C3464 DVDD a_n71_n1840# 0.192782f
C3465 a_n71_n600# a_n71_n1840# 0.001197f
C3466 a_2995_n4294# a_2363_n2734# 3.12e-19
C3467 a_5456_n3308# A8 3.08e-21
C3468 B7 B11 0.001479f
C3469 a_2315_n4255# a_1201_n4294# 0.024621f
C3470 a_6023_n1814# B14 0.056624f
C3471 a_1261_n4320# a_n131_n4294# 0.011053f
C3472 B15 a_3736_n828# 3.18e-19
C3473 a_1968_n4294# a_1201_n3054# 1.81e-21
C3474 a_1467_n3674# a_2995_n4294# 3.6e-21
C3475 B5 a_1479_n2734# 0.002612f
C3476 a_143_n2276# a_1261_n4320# 1.44e-20
C3477 a_5192_n828# a_3543_n342# 3.51e-20
C3478 DVDD a_4523_n574# 0.005567f
C3479 a_3832_n1194# a_3946_n1066# 2.79e-19
C3480 a_4000_n1194# a_3874_n1220# 0.045338f
C3481 a_1997_n1194# a_2273_n254# 0.001323f
C3482 a_636_n3054# a_2254_n1194# 1.34e-20
C3483 B9 a_3655_n1516# 1.39e-19
C3484 A11 a_4523_n3054# 3.39e-19
C3485 DVDD a_6023_n1494# 5.73e-19
C3486 a_143_n2276# B15 9.21e-20
C3487 DVDD a_1557_n2434# 0.369711f
C3488 a_4000_n1194# a_3946_174# 7.6e-20
C3489 a_541_n2434# a_101_n3674# 1.67e-20
C3490 a_2459_n2734# a_1201_n3054# 0.009339f
C3491 B11 a_5402_n3546# 7.19e-19
C3492 a_2363_n2734# a_1201_n4294# 1.46e-22
C3493 a_2273_n2734# a_n131_n4294# 0.034838f
C3494 a_5819_n2068# a_3543_n342# 0.003904f
C3495 a_11_n2434# a_n131_n1814# 1.2e-19
C3496 a_143_n2276# a_2273_n2734# 0.058245f
C3497 B13 a_3874_n1220# 1.11e-19
C3498 a_2995_n4294# a_2350_n2434# 1.39e-19
C3499 a_2254_n2434# a_1968_n1814# 4.57e-19
C3500 DVDD a_1997_46# 8.16e-19
C3501 a_1467_n3674# a_1201_n4294# 9.84e-21
C3502 a_966_n3674# a_n131_n4294# 1.65e-19
C3503 a_2995_n4294# B5 0.005611f
C3504 a_2995_n4294# a_4000_n828# 6.25e-19
C3505 a_4204_n3054# a_6023_n4294# 1.35e-19
C3506 a_541_46# a_894_46# 2.18e-19
C3507 a_1968_n4294# a_636_n4294# 1.72e-19
C3508 A12 a_3874_20# 0.021138f
C3509 B13 a_3946_174# 0.17279f
C3510 A13 a_636_n574# 2.02e-20
C3511 DVDD a_4697_412# 5e-19
C3512 a_5456_46# a_5360_46# 0.023012f
C3513 Cin a_3904_46# 1.26e-19
C3514 a_5402_n3546# a_4204_n3054# 0.219575f
C3515 a_2273_n2734# a_1641_n3308# 0.001272f
C3516 a_5192_n3674# a_3543_n2822# 1.65e-19
C3517 a_4697_n3674# a_3669_n2822# 9.84e-21
C3518 a_3322_n1582# a_4363_n828# 0.001272f
C3519 a_3765_n3080# a_3543_n342# 6.14e-21
C3520 a_3669_n2822# a_3669_n342# 2.45e-20
C3521 a_4204_n574# a_4000_n828# 5.14e-19
C3522 a_3861_n3080# a_2908_n600# 4.82e-21
C3523 a_3368_n1448# a_2995_n4294# 3.4e-19
C3524 a_5360_n2434# a_3946_n2306# 0.031298f
C3525 B14 a_5288_n828# 2.91e-19
C3526 B13 a_4523_n574# 0.007771f
C3527 a_3904_46# a_3669_n342# 3.97e-19
C3528 a_n131_n574# a_1201_n1814# 0.006573f
C3529 B5 a_1201_n4294# 6.28e-19
C3530 a_101_n1194# a_n131_n574# 2.05e-19
C3531 a_636_n1814# a_1261_n600# 5.78e-19
C3532 a_5456_n3308# a_4204_n3054# 0.087066f
C3533 a_1641_n3674# a_636_n4294# 0.033252f
C3534 a_1997_n3674# a_101_n3674# 5.42e-21
C3535 DVDD A15 0.480085f
C3536 B3 a_1261_n600# 7.54e-19
C3537 a_2273_n254# a_3861_n600# 1.64e-19
C3538 a_636_n3054# a_1647_n3054# 2.35e-19
C3539 A14 a_5819_n1194# 0.050725f
C3540 A7 a_2995_n4294# 0.006765f
C3541 a_966_n2068# a_n131_n1814# 4.28e-20
C3542 DVDD a_5819_n828# 0.162119f
C3543 DVDD B8 0.775697f
C3544 a_101_46# a_185_46# 0.067562f
C3545 a_3874_n2460# a_3669_n2822# 7.1e-20
C3546 a_3946_n2306# a_3543_n2822# 7.63e-19
C3547 a_143_n2276# a_3177_n1814# 0.087128f
C3548 a_894_n2434# B4 7.33e-20
C3549 a_966_n2434# a_101_n2434# 3.46e-19
C3550 a_894_n2434# a_636_n3054# 2.34e-19
C3551 Cin a_2363_n254# 8.07e-19
C3552 a_4204_n574# a_5456_46# 7.7e-21
C3553 a_1557_46# a_2908_n600# 2.26e-20
C3554 B9 a_5773_n3054# 3.52e-21
C3555 a_101_46# a_11_412# 0.006823f
C3556 A9 a_3669_n342# 1.38e-19
C3557 a_2273_n2734# a_1968_n1814# 4.1e-20
C3558 a_1261_n600# a_1291_n574# 0.025037f
C3559 a_2790_n3928# a_2995_n4294# 0.001141f
C3560 a_2254_n3674# a_1557_n3674# 0.051953f
C3561 A14 a_3322_n1582# 5.21e-20
C3562 a_3322_n1582# a_3543_n2822# 3.04e-20
C3563 B9 a_4363_n2068# 0.020016f
C3564 A7 a_1201_n4294# 0.077871f
C3565 DVDD a_1997_n3308# 0.154852f
C3566 DVDD a_1997_n1194# 8.16e-19
C3567 A5 a_1557_n3674# 2.88e-19
C3568 a_4204_n3054# a_5288_n3308# 2.9e-19
C3569 a_11_n2434# A4 4.78e-19
C3570 a_4000_n1194# A15 0.046632f
C3571 a_3669_n2822# a_n131_n3054# 6.1e-20
C3572 a_3543_n2822# a_1201_n3054# 3.23e-20
C3573 a_3946_n1066# a_4363_n828# 0.030161f
C3574 a_3874_n1220# a_4697_n828# 7.45e-20
C3575 A10 a_3874_n3700# 0.020957f
C3576 B15 a_4523_n1814# 0.007771f
C3577 a_3434_n1546# a_4441_n1814# 0.053796f
C3578 DVDD A10 0.485225f
C3579 a_3874_n2460# A9 0.512147f
C3580 a_2569_n3928# a_n131_n4294# 0.001075f
C3581 a_143_n2276# a_2569_n3928# 0.003803f
C3582 a_636_n574# a_2350_412# 1.35e-20
C3583 A13 B15 0.004004f
C3584 B13 A15 0.007762f
C3585 a_1997_n3674# a_1557_n2434# 7.6e-20
C3586 B5 a_2315_n1775# 1.39e-19
C3587 a_2273_n254# a_1201_n4294# 1.12e-20
C3588 a_143_n2276# a_143_n1036# 0.003981f
C3589 a_1647_n1814# a_2273_n254# 3.9e-20
C3590 a_2254_n2434# a_2350_n2068# 0.004869f
C3591 a_1997_n2068# a_2422_n2068# 1.31e-19
C3592 Cin a_2350_n828# 7.72e-21
C3593 B14 a_3543_n342# 0.057188f
C3594 a_541_n1194# a_894_n1194# 2.18e-19
C3595 a_4691_n1814# a_4441_n1814# 0.025037f
C3596 A2 a_n41_n574# 7.55e-19
C3597 a_5402_n1066# a_5456_46# 1.67e-20
C3598 a_4691_n3054# a_4441_n3054# 0.025037f
C3599 a_636_n4294# a_3543_n2822# 1.07e-20
C3600 B6 a_1557_n3674# 3.07e-19
C3601 A12 a_5773_n1814# 2.8e-21
C3602 a_5855_n3054# a_3861_n3080# 0.00528f
C3603 a_6153_n2068# A8 5.12e-20
C3604 a_2422_n2068# A5 1.05e-19
C3605 a_n131_n4294# a_2569_n1775# 2.63e-20
C3606 A1 a_2273_n254# 4.12e-19
C3607 B0 a_1201_n574# 4.3e-20
C3608 a_3177_n1814# a_1968_n1814# 1.52e-19
C3609 a_143_n2276# a_2569_n1775# 0.104916f
C3610 a_5192_n3674# a_3946_n3546# 3.2e-20
C3611 a_5288_n3674# a_3874_n3700# 2.34e-19
C3612 a_966_n2068# A4 1.05e-19
C3613 a_4000_n3674# a_3669_n2822# 0.001261f
C3614 a_1557_n3674# a_143_n3516# 0.005791f
C3615 a_3946_n1066# A14 0.001406f
C3616 a_n41_n4294# a_636_n4294# 1.77e-19
C3617 a_541_n1194# a_143_n1036# 0.045338f
C3618 DVDD a_3861_n600# 1.67723f
C3619 a_3904_n3674# a_4000_n3308# 0.02283f
C3620 B14 a_5288_n1194# 7.33e-20
C3621 a_2422_46# a_2254_46# 0.00792f
C3622 a_3322_n4062# B10 2.25e-20
C3623 a_5360_n3674# a_5192_n3674# 0.00792f
C3624 DVDD a_541_n3674# 0.002071f
C3625 DVDD a_5360_46# 0.234826f
C3626 a_5819_n3308# a_3543_n342# 2.31e-19
C3627 a_2995_n4294# a_4691_n4294# 2.91e-20
C3628 a_798_n1194# a_n131_n1814# 0.001991f
C3629 A3 a_2908_n600# 5.91e-19
C3630 a_3434_n1546# a_3322_n4062# 4.1e-20
C3631 A8 a_3861_n3080# 0.025968f
C3632 a_3874_20# a_4000_412# 0.112124f
C3633 a_3946_174# a_3904_46# 0.055111f
C3634 a_2254_n2434# a_2315_n4255# 7.07e-21
C3635 a_1479_n254# a_143_n1036# 5.41e-19
C3636 a_2254_n3674# a_1968_n4294# 1.54e-19
C3637 B9 a_2908_n600# 8.43e-21
C3638 A2 a_966_n1194# 7.66e-19
C3639 a_3946_n2306# a_3946_n3546# 0.007318f
C3640 a_3874_n2460# a_5402_n3546# 1.11e-19
C3641 a_2995_n4294# a_3874_n3700# 0.008003f
C3642 a_4441_n1814# a_4441_n3054# 0.002078f
C3643 a_5773_n1814# a_3861_n3080# 1.74e-20
C3644 a_4204_n3054# a_4000_n2434# 7.87e-20
C3645 B1 a_143_n2276# 0.001432f
C3646 B7 a_n131_n3054# 8.88e-19
C3647 DVDD a_2995_n4294# 1.93905f
C3648 a_636_n1814# a_1557_46# 0.002601f
C3649 a_3736_n1194# B15 6.11e-20
C3650 a_143_n1036# a_1968_n1814# 8.25e-20
C3651 Cin a_2569_n1448# 0.003803f
C3652 a_2273_n254# a_2315_n1775# 0.236061f
C3653 a_2350_n2068# a_2273_n2734# 1.21e-20
C3654 B3 a_1557_46# 4.05e-20
C3655 a_3711_n254# a_1201_n574# 9.58e-21
C3656 a_2422_n3308# a_2273_n2734# 1.91e-19
C3657 A2 a_2273_n254# 5.21e-20
C3658 a_143_n1036# a_966_412# 2.91e-20
C3659 DVDD a_4204_n574# 0.781074f
C3660 a_143_n2276# a_1641_n828# 9.97e-19
C3661 B11 a_4441_n4294# 0.2191f
C3662 a_143_n3516# a_315_n3054# 8.43e-19
C3663 a_3874_n3700# a_1201_n4294# 8.93e-21
C3664 a_1557_n3674# a_n131_n4294# 0.002594f
C3665 a_315_n1814# a_n131_n1814# 0.003681f
C3666 a_5456_n828# a_5192_n828# 1.31e-19
C3667 a_143_n2276# a_1557_n3674# 0.001513f
C3668 B11 a_3861_n3080# 8.88e-19
C3669 B13 a_3861_n600# 0.033034f
C3670 a_1968_n1814# a_2569_n1775# 0.190276f
C3671 a_n71_n4320# a_1968_n4294# 1.26e-20
C3672 DVDD a_1201_n4294# 0.367021f
C3673 A12 a_5360_n1194# 2.18e-20
C3674 DVDD a_1647_n1814# 0.008551f
C3675 a_636_n574# a_n41_n574# 4.33e-19
C3676 B7 a_101_n3674# 7.19e-19
C3677 B13 a_5360_46# 2.55e-19
C3678 a_5192_n2434# a_5456_n2434# 8.12e-20
C3679 a_3711_n2734# a_3322_n4062# 7.42e-19
C3680 a_798_n2434# B4 0.078639f
C3681 a_3736_n2068# a_2995_n4294# 4.55e-19
C3682 A1 a_1997_n828# 8.69e-21
C3683 a_3832_n2068# a_3946_n2306# 4.35e-21
C3684 a_894_n2068# a_101_n2434# 4.35e-21
C3685 a_798_n2434# a_636_n3054# 0.012687f
C3686 A4 a_n131_n1814# 0.012262f
C3687 B6 a_1968_n4294# 1.57e-20
C3688 a_3832_n3308# a_2995_n4294# 7.4e-20
C3689 a_4000_n1194# a_2995_n4294# 9.16e-19
C3690 a_2254_n2434# a_2350_n2434# 0.005587f
C3691 a_3736_46# a_4000_46# 8.12e-20
C3692 a_4441_n4294# a_4204_n3054# 5.74e-19
C3693 a_1557_n3674# a_1641_n3308# 0.030161f
C3694 a_5456_n2068# B8 0.017703f
C3695 B1 a_1479_n254# 0.002612f
C3696 a_2254_n2434# B5 0.077428f
C3697 DVDD A1 0.443246f
C3698 A1 a_n71_n600# 1.38e-21
C3699 Cin a_1261_n600# 9.92e-19
C3700 A0 Cin 0.472133f
C3701 a_1291_n1814# A3 0.007493f
C3702 a_4000_412# a_4363_412# 0.009846f
C3703 a_3861_n3080# a_4204_n3054# 0.182595f
C3704 a_4441_n3054# a_3322_n4062# 6.57e-19
C3705 a_2995_n4294# a_1291_n3054# 2.18e-19
C3706 a_2315_n4255# a_2273_n2734# 0.236061f
C3707 a_1968_n4294# a_143_n3516# 8.25e-20
C3708 A5 a_2422_n2434# 7.66e-19
C3709 a_2995_n4294# a_4697_n3308# 1.06e-20
C3710 a_185_n3308# a_n131_n1814# 2.31e-19
C3711 B2 a_143_n2276# 7.65e-19
C3712 DVDD a_1467_n3308# 4.94e-19
C3713 B13 a_2995_n4294# 3.1e-19
C3714 a_1557_n2434# A9 2.18e-20
C3715 a_4000_n1194# a_4204_n574# 4.76e-20
C3716 DVDD a_185_n1194# 0.003788f
C3717 a_1201_n574# a_2908_n600# 2.14e-19
C3718 a_1201_n1814# a_n131_n1814# 1.11131f
C3719 a_n131_n574# a_3543_n342# 8.62e-20
C3720 a_101_n1194# a_n131_n1814# 0.034089f
C3721 a_798_n1194# A4 1.29e-20
C3722 a_2422_n2068# a_143_n2276# 3.86e-19
C3723 a_3946_n1066# a_2254_n1194# 2.97e-20
C3724 a_541_412# a_798_46# 0.02283f
C3725 a_143_n1036# a_1467_n828# 5.15e-20
C3726 a_4000_n3674# a_5402_n3546# 5.42e-21
C3727 a_4363_n3674# a_3946_n3546# 0.06777f
C3728 A14 a_6153_n828# 5.12e-20
C3729 A15 a_3904_46# 1.29e-20
C3730 a_2273_n2734# a_2363_n2734# 0.010797f
C3731 B13 a_4204_n574# 0.046267f
C3732 DVDD a_5402_n1066# 0.389179f
C3733 B14 a_6153_n1194# 3.15e-19
C3734 Cin a_3226_n1582# 0.00255f
C3735 a_1291_n3054# a_1201_n4294# 2.26e-19
C3736 a_798_n2434# A6 1.29e-20
C3737 a_1647_n3054# a_1201_n3054# 0.001897f
C3738 a_315_n3054# a_n131_n4294# 2.52e-19
C3739 a_1641_n3674# a_143_n3516# 9.15e-19
C3740 a_5402_174# a_5456_412# 0.004108f
C3741 a_n41_n1814# a_n71_n3080# 3.47e-20
C3742 a_2569_n4255# a_2995_n4294# 0.096027f
C3743 B2 a_541_n1194# 0.005557f
C3744 a_3543_n342# B10 2.66e-19
C3745 A7 a_2254_n2434# 1.29e-20
C3746 a_1261_n4320# B5 3.66e-21
C3747 a_798_n1194# a_101_n1194# 0.057934f
C3748 a_636_n1814# A3 0.51166f
C3749 a_3434_n1546# a_3543_n342# 0.031799f
C3750 a_3226_n1582# a_3669_n342# 1.29e-20
C3751 a_3655_n1516# a_2908_n600# 6.53e-19
C3752 a_636_n574# a_2273_n254# 3.49e-19
C3753 a_2254_n3674# a_3543_n2822# 1.02e-19
C3754 A3 B3 1.25275f
C3755 DVDD a_2315_n1775# 0.194591f
C3756 a_1997_n1194# a_1641_n1194# 0.008475f
C3757 B7 a_1557_n2434# 4.05e-20
C3758 A7 a_3904_n3674# 9.68e-20
C3759 a_4363_46# a_4000_46# 0.008475f
C3760 A1 B13 2.72e-20
C3761 B1 A13 2.72e-20
C3762 DVDD A2 0.513733f
C3763 A2 a_n71_n600# 0.001913f
C3764 a_2273_n2734# a_2350_n2434# 6.08e-20
C3765 A15 A9 0.001672f
C3766 a_2569_n4255# a_1201_n4294# 1.29e-20
C3767 B15 a_4000_n828# 0.005326f
C3768 a_1968_n4294# a_n131_n4294# 0.031799f
C3769 a_1997_n3674# a_2995_n4294# 8.26e-19
C3770 a_143_n2276# a_1968_n4294# 0.299183f
C3771 B5 a_2273_n2734# 0.001085f
C3772 DVDD a_5855_n574# 0.005567f
C3773 a_4691_n1814# a_3543_n342# 0.017157f
C3774 A9 B8 1.74e-19
C3775 B9 A8 2.69e-19
C3776 A10 a_3669_n2822# 1.6e-19
C3777 a_2254_n2434# a_2273_n254# 2.41e-19
C3778 a_4000_n1194# a_5402_n1066# 5.42e-21
C3779 a_2422_n1194# a_2273_n254# 4.57e-19
C3780 A8 a_5192_n2434# 7.66e-19
C3781 A3 a_1291_n574# 7.81e-20
C3782 B2 a_1968_n1814# 1.57e-20
C3783 a_5819_n2434# B10 8.1e-22
C3784 a_315_n1814# a_1201_n1814# 1.83e-19
C3785 DVDD a_3685_n1775# 8.63e-19
C3786 a_n41_n1814# a_636_n1814# 1.77e-19
C3787 A7 a_1261_n4320# 0.084607f
C3788 a_143_n2276# a_2459_n2734# 6.86e-19
C3789 a_3874_n2460# a_4000_n2434# 0.045338f
C3790 a_3946_n2306# a_3832_n2434# 3.53e-19
C3791 A12 a_5773_n574# 0.081598f
C3792 a_2995_n4294# a_3736_n2434# 9.92e-19
C3793 a_2273_n254# a_2350_46# 6.08e-20
C3794 a_1997_n3674# a_1201_n4294# 0.001261f
C3795 A11 a_3736_n3674# 7.66e-19
C3796 A4 a_185_n3308# 7.78e-19
C3797 DVDD a_1467_46# 3.22e-21
C3798 Cin a_541_46# 0.045338f
C3799 B0 a_894_46# 7.33e-20
C3800 a_2995_n4294# a_4697_n828# 8.18e-21
C3801 A0 a_966_46# 7.66e-19
C3802 a_101_n1194# A4 0.003351f
C3803 a_1641_n2434# B3 2.95e-21
C3804 DVDD a_3368_n4255# 0.001765f
C3805 a_1479_n1494# a_1261_n1840# 0.007234f
C3806 a_3832_n828# a_4000_n828# 2.18e-19
C3807 A7 a_2273_n2734# 0.037805f
C3808 a_n41_n4294# a_n71_n4320# 0.025037f
C3809 B11 B9 0.005115f
C3810 a_5456_n3674# a_3543_n2822# 0.001186f
C3811 a_4441_n3054# a_3543_n342# 8.88e-21
C3812 a_3861_n3080# a_3669_n342# 5.47e-21
C3813 a_3322_n1582# a_5192_n828# 1.79e-20
C3814 a_4204_n574# a_4697_n828# 5.15e-20
C3815 a_5456_n2068# a_2995_n4294# 0.091184f
C3816 B6 a_n41_n4294# 0.056624f
C3817 a_5360_n2434# a_5402_n2306# 0.057766f
C3818 A6 a_11_n3308# 5.12e-20
C3819 B14 a_5456_n828# 0.017703f
C3820 a_143_n2276# a_2422_n2434# 7.48e-19
C3821 a_3904_46# a_3861_n600# 3.5e-19
C3822 a_1557_n1194# a_n131_n574# 6.4e-19
C3823 a_101_n1194# a_1201_n1814# 0.003559f
C3824 a_636_n1814# a_1201_n574# 1.04e-19
C3825 a_6153_n3308# a_4204_n3054# 1.23e-20
C3826 a_n41_n4294# a_143_n3516# 1.35e-19
C3827 a_3543_n342# a_4000_n2068# 0.001046f
C3828 B3 a_1201_n574# 0.00216f
C3829 B8 a_5402_n3546# 6.9e-19
C3830 a_5456_n2068# a_4204_n574# 6.58e-21
C3831 a_1641_n2068# a_n131_n1814# 0.001068f
C3832 a_6023_n3054# B10 3.35e-19
C3833 B7 a_1997_n3308# 0.005326f
C3834 Cin a_1557_46# 0.081577f
C3835 a_2273_n254# a_2273_n2734# 6.99e-20
C3836 B9 a_4204_n3054# 0.046267f
C3837 a_4441_n4294# a_3874_n2460# 9.91e-21
C3838 a_3434_n4026# a_2995_n4294# 0.305534f
C3839 DVDD a_11_n1194# 2.33e-19
C3840 DVDD a_636_n574# 0.899769f
C3841 B1 a_2350_412# 2.91e-19
C3842 A0 a_101_46# 0.780011f
C3843 A1 a_2422_412# 1.05e-19
C3844 a_636_n574# a_n71_n600# 0.063303f
C3845 a_101_46# a_1261_n600# 0.005909f
C3846 a_4204_n3054# a_5192_n2434# 1.96e-19
C3847 a_5402_n2306# a_3543_n2822# 2.69e-19
C3848 A0 a_n71_n1840# 2.8e-21
C3849 a_2995_n4294# a_3669_n2822# 0.025086f
C3850 a_3874_n2460# a_3861_n3080# 0.289331f
C3851 A14 a_5402_n2306# 6.58e-20
C3852 a_3946_n2306# a_3765_n3080# 0.076462f
C3853 a_3177_n1814# a_3368_n1448# 2.88e-19
C3854 a_1641_n2434# a_101_n2434# 1.11e-20
C3855 Cin a_2543_n254# 6.47e-19
C3856 a_966_n2434# a_1557_n2434# 3.2e-20
C3857 A2 a_185_46# 4.33e-21
C3858 A11 B11 1.25275f
C3859 a_2350_n1194# a_2254_n1194# 0.005587f
C3860 a_1201_n574# a_1291_n574# 0.074717f
C3861 a_n131_n574# a_1647_n574# 0.005159f
C3862 a_2254_n3674# a_3946_n3546# 2.97e-20
C3863 a_3874_n2460# a_3904_n2434# 0.062548f
C3864 a_3627_n254# a_3543_n342# 2.77e-20
C3865 a_2543_n2734# a_1201_n3054# 3.31e-19
C3866 a_2459_n254# a_3765_n600# 9.58e-21
C3867 A10 a_6023_n4294# 0.007489f
C3868 DVDD a_2254_n2434# 0.247054f
C3869 a_3322_n1582# a_3765_n3080# 4.56e-21
C3870 DVDD a_2350_n3308# 4.94e-19
C3871 DVDD a_11_n828# 5.28e-19
C3872 a_636_n574# a_1467_412# 7.45e-20
C3873 a_3874_n3700# a_3904_n3674# 0.06247f
C3874 a_3543_n2822# a_n131_n4294# 0.011993f
C3875 a_3765_n3080# a_1201_n3054# 0.001811f
C3876 a_3861_n3080# a_n131_n3054# 7.7e-20
C3877 a_3669_n2822# a_1201_n4294# 8.04e-19
C3878 a_143_n2276# a_3543_n2822# 1.59e-19
C3879 a_636_n3054# a_n131_n574# 4.68e-22
C3880 a_143_n2276# a_1467_n1194# 1.36e-20
C3881 DVDD a_3904_n3674# 0.247054f
C3882 A10 a_5402_n3546# 0.780011f
C3883 a_185_n2434# a_n131_n1814# 0.001123f
C3884 A11 a_4204_n3054# 0.011053f
C3885 a_n41_n574# a_143_n1036# 0.002038f
C3886 a_2995_n4294# A9 0.082881f
C3887 a_n41_n4294# a_n131_n4294# 0.096176f
C3888 a_315_n4294# a_1201_n4294# 1.83e-19
C3889 a_541_46# a_966_46# 8.12e-20
C3890 B12 a_3874_20# 0.014043f
C3891 A12 a_3946_174# 0.001406f
C3892 A10 a_5456_n3308# 0.011819f
C3893 a_5456_n2068# a_5402_n1066# 1.79e-19
C3894 a_3177_n1814# a_2273_n254# 8.15e-19
C3895 B13 a_636_n574# 2.79e-20
C3896 a_4523_n3054# a_4204_n3054# 0.003613f
C3897 a_4691_n3054# a_3322_n4062# 5.44e-19
C3898 a_2315_n4255# a_1557_n3674# 0.027489f
C3899 DVDD a_5192_412# 6.81e-19
C3900 A1 a_3904_46# 9.68e-20
C3901 a_3434_n1546# a_4691_n1494# 3.05e-19
C3902 S15 a_2543_n254# 3.11e-20
C3903 a_5773_n4294# a_6023_n3054# 3.47e-20
C3904 a_5855_n1814# a_5773_n1814# 0.006406f
C3905 DVDD a_1261_n4320# 0.184562f
C3906 a_143_n2276# a_185_n2068# 0.091046f
C3907 a_5855_n3054# a_5773_n3054# 0.006406f
C3908 a_n131_n1814# a_3543_n342# 0.006998f
C3909 a_3322_n1582# a_3736_46# 2.27e-20
C3910 a_3589_n1448# a_1968_n1814# 3.16e-20
C3911 a_3736_n3308# a_4000_n3308# 1.31e-19
C3912 a_3832_n3308# a_3904_n3674# 0.004869f
C3913 a_5288_n3674# a_5402_n3546# 3.78e-19
C3914 a_3874_n3700# a_2273_n2734# 7.5e-21
C3915 a_3946_n1066# a_3765_n3080# -5.88e-38
C3916 a_1291_n4294# a_636_n4294# 6.24e-19
C3917 DVDD B15 0.619467f
C3918 DVDD a_5819_n3674# 0.001386f
C3919 Cin A3 0.001563f
C3920 A5 a_1647_n3054# 1.5e-19
C3921 a_966_n1194# a_143_n1036# 1.32e-19
C3922 B14 a_5819_n1194# 0.021045f
C3923 B7 a_2995_n4294# 0.004799f
C3924 a_4000_n3308# a_4363_n3308# 0.009846f
C3925 a_1467_n3674# a_1557_n3674# 0.006958f
C3926 DVDD a_2273_n2734# 1.15045f
C3927 a_1557_46# a_966_46# 3.2e-20
C3928 A13 a_4363_n828# 1.58e-21
C3929 a_5360_n3674# a_5456_n3674# 0.023012f
C3930 a_3669_n342# a_4363_n1194# 9.33e-19
C3931 a_101_46# a_541_46# 0.044963f
C3932 DVDD a_966_n3674# 9.02e-20
C3933 A3 a_3669_n342# 7.21e-20
C3934 a_3874_n1220# a_3904_n2434# 1.17e-20
C3935 a_4204_n574# a_5819_46# 1.55e-21
C3936 A8 a_5773_n3054# 0.081598f
C3937 a_143_n1036# a_2273_n254# 0.01799f
C3938 a_11_n2434# B4 3.15e-19
C3939 B9 a_3669_n342# 2.37e-19
C3940 a_5773_n1814# a_5773_n3054# 0.001197f
C3941 a_1641_412# a_1997_412# 0.009846f
C3942 B14 a_3322_n1582# 2.25e-20
C3943 B7 a_1201_n4294# 0.081283f
C3944 A14 a_6023_n574# 7.55e-19
C3945 a_1261_n4320# a_1291_n3054# 9.75e-20
C3946 DVDD a_11_n2068# 5.28e-19
C3947 B5 a_1557_n3674# 3.5e-19
C3948 a_185_n2434# A4 0.050725f
C3949 a_4000_n1194# B15 0.005557f
C3950 a_2273_n254# a_2569_n1775# 0.318695f
C3951 a_3874_n2460# a_4363_n1194# 1.55e-21
C3952 a_5456_n3308# a_2995_n4294# 6.58e-21
C3953 a_5360_n3674# a_5402_n2306# 1.16e-19
C3954 DVDD a_3832_n828# 4.94e-19
C3955 a_1557_46# a_3946_174# 0.001288f
C3956 a_541_n2068# A2 3.08e-21
C3957 a_n131_n1814# a_1261_n3080# 8.88e-21
C3958 a_101_n1194# a_798_46# 9.75e-22
C3959 a_101_46# a_1557_46# 0.003292f
C3960 a_143_n2276# a_2254_n1194# 0.004198f
C3961 a_3874_n2460# B9 1.25937f
C3962 a_2273_n2734# a_1291_n3054# 5.44e-19
C3963 a_143_n3516# a_1647_n3054# 0.003613f
C3964 a_3946_n3546# a_n131_n4294# 1.19e-20
C3965 a_143_n2276# a_3946_n3546# 1.42e-20
C3966 B7 a_1467_n3308# 4.23e-20
C3967 B13 B15 0.005115f
C3968 a_3946_n2306# a_4697_n2434# 0.006958f
C3969 a_3874_n2460# a_5192_n2434# 3.15e-19
C3970 A11 a_4697_n3674# 5.03e-19
C3971 a_2315_n4255# a_1968_n4294# 0.153192f
C3972 A12 a_5819_n828# 7.78e-19
C3973 DVDD a_3177_n1814# 0.145407f
C3974 a_1557_n2434# a_3904_n2434# 2.97e-20
C3975 a_894_n2434# a_143_n3516# 1.66e-19
C3976 a_966_n2068# B4 3.18e-19
C3977 a_3543_n2822# a_3685_n4255# 9.8e-19
C3978 A3 a_n131_n3054# 1.7e-21
C3979 B12 a_5773_n1814# 8.21e-21
C3980 B2 a_n41_n574# 3.35e-19
C3981 A7 a_1557_n3674# 0.791917f
C3982 a_2422_n2068# B5 3.18e-19
C3983 B1 a_2273_n254# 0.001085f
C3984 Cin a_1201_n574# 0.006883f
C3985 a_5773_n3054# a_4204_n3054# 0.001762f
C3986 a_2569_n4255# a_2273_n2734# 0.318695f
C3987 B10 DGND 0.973708f
C3988 A10 DGND 0.991087f
C3989 B11 DGND 0.870336f
C3990 A11 DGND 1.01949f
C3991 B7 DGND 0.870336f
C3992 A7 DGND 1.01949f
C3993 B6 DGND 0.973999f
C3994 A6 DGND 0.991699f
C3995 B8 DGND 0.98773f
C3996 A8 DGND 1.04702f
C3997 B9 DGND 0.824151f
C3998 A9 DGND 0.977237f
C3999 B5 DGND 0.824468f
C4000 A5 DGND 0.977254f
C4001 B4 DGND 0.994934f
C4002 A4 DGND 1.03251f
C4003 B14 DGND 0.979861f
C4004 A14 DGND 1.0418f
C4005 B15 DGND 0.852393f
C4006 A15 DGND 1.00441f
C4007 B3 DGND 0.852117f
C4008 A3 DGND 1.00406f
C4009 B2 DGND 0.978379f
C4010 A2 DGND 1.02466f
C4011 S15 DGND 0.143153f
C4012 B12 DGND 0.987081f
C4013 A12 DGND 0.998982f
C4014 B13 DGND 0.855886f
C4015 A13 DGND 1.00181f
C4016 B1 DGND 0.855934f
C4017 A1 DGND 1.00179f
C4018 Cin DGND 1.39034f
C4019 B0 DGND 0.987659f
C4020 A0 DGND 0.998637f
C4021 DVDD DGND 60.932087f
C4022 a_6023_n4294# DGND 0.004578f
C4023 a_5855_n4294# DGND 0.001767f
C4024 a_4691_n4294# DGND 0.003702f
C4025 a_4523_n4294# DGND 0.001767f
C4026 a_3685_n4255# DGND 2.7e-19
C4027 a_3368_n4255# DGND 6.44e-19
C4028 a_6023_n3974# DGND 0.005523f
C4029 a_4691_n3974# DGND 0.005523f
C4030 a_2783_n4255# DGND 6.44e-19
C4031 a_2497_n4255# DGND 2.7e-19
C4032 a_3589_n3928# DGND 0.003343f
C4033 a_3368_n3928# DGND 0.003279f
C4034 a_1647_n4294# DGND 0.001767f
C4035 a_1291_n4294# DGND 0.003702f
C4036 a_315_n4294# DGND 0.001767f
C4037 a_n41_n4294# DGND 0.004578f
C4038 a_2790_n3928# DGND 0.003279f
C4039 a_2569_n3928# DGND 0.003343f
C4040 a_1479_n3974# DGND 0.005523f
C4041 a_147_n3974# DGND 0.005523f
C4042 a_5773_n4294# DGND 0.364177f
C4043 a_4441_n4294# DGND 0.354376f
C4044 a_3655_n3996# DGND 0.303354f
C4045 a_3434_n4026# DGND 0.681093f
C4046 a_3226_n4062# DGND 0.282084f
C4047 a_2569_n4255# DGND 0.282084f
C4048 a_1968_n4294# DGND 0.681093f
C4049 a_2315_n4255# DGND 0.303354f
C4050 a_1261_n4320# DGND 0.354376f
C4051 a_n71_n4320# DGND 0.363945f
C4052 a_6153_n3674# DGND 0.002125f
C4053 a_5819_n3674# DGND 0.159242f
C4054 a_5456_n3674# DGND 0.165381f
C4055 a_5288_n3674# DGND 0.001155f
C4056 a_5192_n3674# DGND 0.002255f
C4057 a_4697_n3674# DGND 0.002142f
C4058 a_4363_n3674# DGND 0.159436f
C4059 a_4000_n3674# DGND 0.163641f
C4060 a_3832_n3674# DGND 8.87e-19
C4061 a_3736_n3674# DGND 0.001946f
C4062 a_2422_n3674# DGND 0.001946f
C4063 a_2350_n3674# DGND 8.87e-19
C4064 a_1997_n3674# DGND 0.163641f
C4065 a_1641_n3674# DGND 0.159436f
C4066 a_1467_n3674# DGND 0.002142f
C4067 a_966_n3674# DGND 0.002255f
C4068 a_894_n3674# DGND 0.001156f
C4069 a_541_n3674# DGND 0.165382f
C4070 a_185_n3674# DGND 0.159097f
C4071 a_11_n3674# DGND 0.002194f
C4072 a_5819_n3308# DGND 0.005381f
C4073 a_5456_n3308# DGND 0.008579f
C4074 a_5360_n3674# DGND 0.239621f
C4075 a_5288_n3308# DGND 1.65e-19
C4076 a_5192_n3308# DGND 1.75e-19
C4077 a_4697_n3308# DGND 2.89e-20
C4078 a_4363_n3308# DGND 0.005269f
C4079 a_4000_n3308# DGND 0.005799f
C4080 a_3904_n3674# DGND 0.23617f
C4081 a_3832_n3308# DGND 2.42e-20
C4082 a_3736_n3308# DGND 2.94e-20
C4083 a_2422_n3308# DGND 2.94e-20
C4084 a_2350_n3308# DGND 2.42e-20
C4085 a_2254_n3674# DGND 0.23617f
C4086 a_1997_n3308# DGND 0.005799f
C4087 a_1641_n3308# DGND 0.005269f
C4088 a_1467_n3308# DGND 2.89e-20
C4089 a_966_n3308# DGND 1.75e-19
C4090 a_894_n3308# DGND 1.66e-19
C4091 a_798_n3674# DGND 0.239626f
C4092 a_541_n3308# DGND 0.008581f
C4093 a_185_n3308# DGND 0.005145f
C4094 a_11_n3308# DGND 1.03e-20
C4095 a_5402_n3546# DGND 1.06588f
C4096 a_3946_n3546# DGND 0.947829f
C4097 a_3874_n3700# DGND 0.974632f
C4098 a_1557_n3674# DGND 0.947829f
C4099 a_636_n4294# DGND 0.974641f
C4100 a_101_n3674# DGND 1.06764f
C4101 a_6023_n3054# DGND 0.00426f
C4102 a_5855_n3054# DGND 0.002829f
C4103 a_4691_n3054# DGND 0.005761f
C4104 a_4523_n3054# DGND 7.64e-19
C4105 a_1647_n3054# DGND 7.64e-19
C4106 a_1291_n3054# DGND 0.005761f
C4107 a_315_n3054# DGND 0.001884f
C4108 a_n41_n3054# DGND 0.005072f
C4109 a_6023_n2734# DGND 0.005804f
C4110 a_4691_n2734# DGND 0.00572f
C4111 a_4204_n3054# DGND 0.69379f
C4112 a_3322_n4062# DGND 0.534062f
C4113 a_3795_n2734# DGND 0.003554f
C4114 a_3711_n2734# DGND 0.001843f
C4115 a_3627_n2734# DGND 0.003255f
C4116 a_2543_n2734# DGND 0.003255f
C4117 a_2459_n2734# DGND 0.001843f
C4118 a_2363_n2734# DGND 0.003554f
C4119 a_2273_n2734# DGND 0.534062f
C4120 a_143_n3516# DGND 0.693676f
C4121 a_1479_n2734# DGND 0.00572f
C4122 a_147_n2734# DGND 0.005804f
C4123 a_5773_n3054# DGND 0.362012f
C4124 a_4441_n3054# DGND 0.329488f
C4125 a_3861_n3080# DGND 0.48244f
C4126 a_3765_n3080# DGND 0.840461f
C4127 a_3669_n2822# DGND 0.580488f
C4128 a_3543_n2822# DGND 1.12816f
C4129 a_n131_n4294# DGND 1.12851f
C4130 a_1201_n4294# DGND 0.580488f
C4131 a_1201_n3054# DGND 0.840461f
C4132 a_n131_n3054# DGND 0.483618f
C4133 a_1261_n3080# DGND 0.329488f
C4134 a_n71_n3080# DGND 0.361766f
C4135 a_6153_n2434# DGND 0.002125f
C4136 a_5819_n2434# DGND 0.164229f
C4137 a_5456_n2434# DGND 0.16997f
C4138 a_5288_n2434# DGND 0.001261f
C4139 a_5192_n2434# DGND 0.002341f
C4140 a_4697_n2434# DGND 0.00213f
C4141 a_4363_n2434# DGND 0.158265f
C4142 a_4000_n2434# DGND 0.162762f
C4143 a_3832_n2434# DGND 8.34e-19
C4144 a_3736_n2434# DGND 0.001875f
C4145 a_2422_n2434# DGND 0.001875f
C4146 a_2350_n2434# DGND 8.34e-19
C4147 a_1997_n2434# DGND 0.162839f
C4148 a_1641_n2434# DGND 0.158297f
C4149 a_1467_n2434# DGND 0.002131f
C4150 a_966_n2434# DGND 0.002355f
C4151 a_894_n2434# DGND 0.001274f
C4152 a_541_n2434# DGND 0.17035f
C4153 a_185_n2434# DGND 0.162453f
C4154 a_11_n2434# DGND 0.002316f
C4155 a_5819_n2068# DGND 0.010649f
C4156 a_5456_n2068# DGND 0.012447f
C4157 a_5360_n2434# DGND 0.234031f
C4158 a_5288_n2068# DGND 2.85e-20
C4159 a_5192_n2068# DGND 4.22e-20
C4160 a_4697_n2068# DGND 9.63e-21
C4161 a_4363_n2068# DGND 0.003634f
C4162 a_4000_n2068# DGND 0.004836f
C4163 a_3904_n2434# DGND 0.234352f
C4164 a_2254_n2434# DGND 0.234352f
C4165 a_1997_n2068# DGND 0.004843f
C4166 a_1641_n2068# DGND 0.003555f
C4167 a_966_n2068# DGND 9.21e-20
C4168 a_894_n2068# DGND 9.13e-20
C4169 a_798_n2434# DGND 0.234749f
C4170 a_541_n2068# DGND 0.012812f
C4171 a_185_n2068# DGND 0.009299f
C4172 a_11_n2068# DGND 2.84e-20
C4173 a_5402_n2306# DGND 1.14907f
C4174 a_2995_n4294# DGND 2.50689f
C4175 a_3946_n2306# DGND 0.94105f
C4176 a_3874_n2460# DGND 0.926267f
C4177 a_1557_n2434# DGND 0.941071f
C4178 a_636_n3054# DGND 0.926598f
C4179 a_101_n2434# DGND 1.15723f
C4180 a_6023_n1814# DGND 0.006666f
C4181 a_5855_n1814# DGND 0.00452f
C4182 a_4691_n1814# DGND 0.004883f
C4183 a_4523_n1814# DGND 0.00205f
C4184 a_3685_n1775# DGND 2.7e-19
C4185 a_3368_n1775# DGND 6.44e-19
C4186 a_6023_n1494# DGND 0.006278f
C4187 a_4691_n1494# DGND 0.005732f
C4188 a_2783_n1775# DGND 6.44e-19
C4189 a_2497_n1775# DGND 2.7e-19
C4190 a_3589_n1448# DGND 0.003343f
C4191 a_3368_n1448# DGND 0.003279f
C4192 a_3177_n1814# DGND 0.077938f
C4193 a_143_n2276# DGND 1.8629f
C4194 a_1647_n1814# DGND 0.001859f
C4195 a_1291_n1814# DGND 0.004192f
C4196 a_315_n1814# DGND 0.003333f
C4197 a_n41_n1814# DGND 0.009716f
C4198 a_2790_n1448# DGND 0.003279f
C4199 a_2569_n1448# DGND 0.003343f
C4200 a_1479_n1494# DGND 0.005748f
C4201 a_147_n1494# DGND 0.006252f
C4202 a_5773_n1814# DGND 0.372814f
C4203 a_4441_n1814# DGND 0.348221f
C4204 a_3655_n1516# DGND 0.296869f
C4205 a_3434_n1546# DGND 0.676995f
C4206 a_3226_n1582# DGND 0.279782f
C4207 a_2569_n1775# DGND 0.278595f
C4208 a_1968_n1814# DGND 0.677066f
C4209 a_2315_n1775# DGND 0.296869f
C4210 a_1261_n1840# DGND 0.347786f
C4211 a_n71_n1840# DGND 0.375866f
C4212 a_6153_n1194# DGND 0.002125f
C4213 a_5819_n1194# DGND 0.160643f
C4214 a_5456_n1194# DGND 0.168023f
C4215 a_5288_n1194# DGND 0.001329f
C4216 a_5192_n1194# DGND 0.002457f
C4217 a_4697_n1194# DGND 0.002142f
C4218 a_4363_n1194# DGND 0.159436f
C4219 a_4000_n1194# DGND 0.163641f
C4220 a_3832_n1194# DGND 8.87e-19
C4221 a_3736_n1194# DGND 0.001946f
C4222 a_2422_n1194# DGND 0.001946f
C4223 a_2350_n1194# DGND 8.87e-19
C4224 a_1997_n1194# DGND 0.163641f
C4225 a_1641_n1194# DGND 0.159436f
C4226 a_1467_n1194# DGND 0.002142f
C4227 a_966_n1194# DGND 0.002457f
C4228 a_894_n1194# DGND 0.001329f
C4229 a_541_n1194# DGND 0.168023f
C4230 a_185_n1194# DGND 0.159964f
C4231 a_11_n1194# DGND 0.002194f
C4232 a_5819_n828# DGND 0.005877f
C4233 a_5456_n828# DGND 0.009535f
C4234 a_5360_n1194# DGND 0.245234f
C4235 a_5288_n828# DGND 1.92e-19
C4236 a_5192_n828# DGND 2e-19
C4237 a_4697_n828# DGND 2.89e-20
C4238 a_4363_n828# DGND 0.005269f
C4239 a_4000_n828# DGND 0.005799f
C4240 a_3832_n828# DGND 2.42e-20
C4241 a_3736_n828# DGND 2.94e-20
C4242 a_2422_n828# DGND 2.94e-20
C4243 a_2350_n828# DGND 2.42e-20
C4244 a_2254_n1194# DGND 0.234325f
C4245 a_1997_n828# DGND 0.005799f
C4246 a_1641_n828# DGND 0.005269f
C4247 a_1467_n828# DGND 2.89e-20
C4248 a_966_n828# DGND 2e-19
C4249 a_894_n828# DGND 1.92e-19
C4250 a_798_n1194# DGND 0.245234f
C4251 a_541_n828# DGND 0.009535f
C4252 a_185_n828# DGND 0.005449f
C4253 a_11_n828# DGND 1.03e-20
C4254 a_5402_n1066# DGND 1.13221f
C4255 a_3946_n1066# DGND 0.935978f
C4256 a_3874_n1220# DGND 1.00335f
C4257 a_1557_n1194# DGND 0.935997f
C4258 a_636_n1814# DGND 1.00563f
C4259 a_101_n1194# DGND 1.13438f
C4260 a_6023_n574# DGND 0.00426f
C4261 a_5855_n574# DGND 0.00242f
C4262 a_4691_n574# DGND 0.005761f
C4263 a_4523_n574# DGND 7.64e-19
C4264 a_1647_n574# DGND 7.64e-19
C4265 a_1291_n574# DGND 0.005761f
C4266 a_315_n574# DGND 0.001854f
C4267 a_n41_n574# DGND 0.005072f
C4268 a_6023_n254# DGND 0.005804f
C4269 a_4691_n254# DGND 0.00572f
C4270 a_4204_n574# DGND 0.693172f
C4271 a_3322_n1582# DGND 0.524285f
C4272 a_3795_n254# DGND 0.003554f
C4273 a_3711_n254# DGND 0.001843f
C4274 a_3627_n254# DGND 0.003262f
C4275 a_2543_n254# DGND 0.003255f
C4276 a_2459_n254# DGND 0.001843f
C4277 a_2363_n254# DGND 0.003554f
C4278 a_2273_n254# DGND 0.52129f
C4279 a_143_n1036# DGND 0.69276f
C4280 a_1479_n254# DGND 0.00572f
C4281 a_147_n254# DGND 0.005804f
C4282 a_5773_n574# DGND 0.359659f
C4283 a_4441_n574# DGND 0.332217f
C4284 a_3861_n600# DGND 0.478399f
C4285 a_3765_n600# DGND 0.840384f
C4286 a_3669_n342# DGND 0.583825f
C4287 a_3543_n342# DGND 0.774217f
C4288 a_2908_n600# DGND 0.680256f
C4289 a_n131_n1814# DGND 0.761377f
C4290 a_1201_n1814# DGND 0.581132f
C4291 a_1201_n574# DGND 0.839838f
C4292 a_n131_n574# DGND 0.477366f
C4293 a_1261_n600# DGND 0.332217f
C4294 a_n71_n600# DGND 0.36066f
C4295 a_6153_46# DGND 0.002125f
C4296 a_5819_46# DGND 0.158063f
C4297 a_5456_46# DGND 0.163195f
C4298 a_5288_46# DGND 8.87e-19
C4299 a_5192_46# DGND 0.001937f
C4300 a_4697_46# DGND 0.002125f
C4301 a_4363_46# DGND 0.15783f
C4302 a_4000_46# DGND 0.162762f
C4303 a_3832_46# DGND 8.34e-19
C4304 a_3736_46# DGND 0.001875f
C4305 a_2422_46# DGND 0.001875f
C4306 a_2350_46# DGND 8.34e-19
C4307 a_1997_46# DGND 0.162762f
C4308 a_1641_46# DGND 0.15783f
C4309 a_1467_46# DGND 0.002125f
C4310 a_966_46# DGND 0.001937f
C4311 a_894_46# DGND 8.87e-19
C4312 a_541_46# DGND 0.163195f
C4313 a_185_46# DGND 0.15797f
C4314 a_11_46# DGND 0.002125f
C4315 a_5819_412# DGND 0.003447f
C4316 a_5456_412# DGND 0.004836f
C4317 a_5360_46# DGND 0.223331f
C4318 a_4363_412# DGND 0.003447f
C4319 a_4000_412# DGND 0.004836f
C4320 a_3904_46# DGND 0.234352f
C4321 a_2254_46# DGND 0.234352f
C4322 a_1997_412# DGND 0.004836f
C4323 a_1641_412# DGND 0.003447f
C4324 a_798_46# DGND 0.223331f
C4325 a_541_412# DGND 0.004836f
C4326 a_185_412# DGND 0.003447f
C4327 a_5402_174# DGND 1.07755f
C4328 a_3946_174# DGND 0.945533f
C4329 a_3874_20# DGND 0.935981f
C4330 a_1557_46# DGND 0.945533f
C4331 a_636_n574# DGND 0.935931f
C4332 a_101_46# DGND 1.07823f
C4333 a_3177_n4294.t0 DGND 0.036409f
C4334 a_3177_n4294.t9 DGND 0.008251f
C4335 a_3177_n4294.t5 DGND 0.02268f
C4336 a_3177_n4294.n0 DGND 0.071595f
C4337 a_3177_n4294.t6 DGND 0.014825f
C4338 a_3177_n4294.t4 DGND 0.010708f
C4339 a_3177_n4294.n1 DGND 0.064557f
C4340 a_3177_n4294.t8 DGND 0.009876f
C4341 a_3177_n4294.t7 DGND 0.015787f
C4342 a_3177_n4294.n2 DGND 0.03061f
C4343 a_3177_n4294.n3 DGND 0.1121f
C4344 a_3177_n4294.t2 DGND 0.00894f
C4345 a_3177_n4294.t3 DGND 0.016664f
C4346 a_3177_n4294.n4 DGND 0.030545f
C4347 a_3177_n4294.n5 DGND 0.034706f
C4348 a_3177_n4294.n6 DGND 2.36783f
C4349 a_3177_n4294.n7 DGND 0.504533f
C4350 a_3177_n4294.t1 DGND 0.039387f
C4351 DVDD.n0 DGND 0.001045f
C4352 DVDD.n1 DGND 0.002178f
C4353 DVDD.n2 DGND 2.23e-19
C4354 DVDD.n3 DGND 0.001172f
C4355 DVDD.t71 DGND 5.49e-19
C4356 DVDD.t431 DGND 1.51e-19
C4357 DVDD.t498 DGND 1.51e-19
C4358 DVDD.n4 DGND 3.12e-19
C4359 DVDD.n5 DGND 0.001184f
C4360 DVDD.n6 DGND 0.001172f
C4361 DVDD.n7 DGND 3.86e-19
C4362 DVDD.n8 DGND 0.001172f
C4363 DVDD.t429 DGND 7.66e-19
C4364 DVDD.n9 DGND 4.15e-19
C4365 DVDD.n10 DGND 0.001172f
C4366 DVDD.t370 DGND 1.51e-19
C4367 DVDD.t422 DGND 1.51e-19
C4368 DVDD.n11 DGND 3.12e-19
C4369 DVDD.t478 DGND 5.49e-19
C4370 DVDD.n12 DGND 0.001052f
C4371 DVDD.n13 DGND 0.001172f
C4372 DVDD.t427 DGND 1.51e-19
C4373 DVDD.t143 DGND 1.51e-19
C4374 DVDD.n14 DGND 3.12e-19
C4375 DVDD.n15 DGND 4.15e-19
C4376 DVDD.n16 DGND 0.00143f
C4377 DVDD.n17 DGND 0.00143f
C4378 DVDD.t34 DGND 7.6e-19
C4379 DVDD.n18 DGND 4.15e-19
C4380 DVDD.n19 DGND 0.001172f
C4381 DVDD.t267 DGND 1.51e-19
C4382 DVDD.t505 DGND 1.51e-19
C4383 DVDD.n20 DGND 3.12e-19
C4384 DVDD.t209 DGND 5.49e-19
C4385 DVDD.n21 DGND 0.001052f
C4386 DVDD.n22 DGND 0.001172f
C4387 DVDD.t36 DGND 1.51e-19
C4388 DVDD.t245 DGND 1.51e-19
C4389 DVDD.n23 DGND 3.12e-19
C4390 DVDD.n24 DGND 4.15e-19
C4391 DVDD.n25 DGND 0.001172f
C4392 DVDD.t175 DGND 7.66e-19
C4393 DVDD.n26 DGND 0.00143f
C4394 DVDD.t9 DGND 7.6e-19
C4395 DVDD.n27 DGND 4.15e-19
C4396 DVDD.n28 DGND 0.001172f
C4397 DVDD.t380 DGND 1.51e-19
C4398 DVDD.t311 DGND 1.51e-19
C4399 DVDD.n29 DGND 3.12e-19
C4400 DVDD.t156 DGND 5.49e-19
C4401 DVDD.n30 DGND 0.001052f
C4402 DVDD.n31 DGND 0.001172f
C4403 DVDD.t161 DGND 1.51e-19
C4404 DVDD.t17 DGND 1.51e-19
C4405 DVDD.n32 DGND 3.12e-19
C4406 DVDD.n33 DGND 4.15e-19
C4407 DVDD.n34 DGND 0.001172f
C4408 DVDD.t309 DGND 7.66e-19
C4409 DVDD.n35 DGND 0.012547f
C4410 DVDD.t471 DGND 7.66e-19
C4411 DVDD.n36 DGND 0.001178f
C4412 DVDD.n37 DGND 3.39e-19
C4413 DVDD.n38 DGND 2.62e-19
C4414 DVDD.n39 DGND 4.15e-19
C4415 DVDD.n40 DGND 4.15e-19
C4416 DVDD.n41 DGND 0.0021f
C4417 DVDD.t293 DGND 0.001258f
C4418 DVDD.n42 DGND 7.9e-19
C4419 DVDD.t395 DGND 3.58e-19
C4420 DVDD.t412 DGND 3.58e-19
C4421 DVDD.n43 DGND 7.77e-19
C4422 DVDD.n44 DGND 0.002427f
C4423 DVDD.t495 DGND 1.51e-19
C4424 DVDD.t330 DGND 1.51e-19
C4425 DVDD.n45 DGND 3.12e-19
C4426 DVDD.n46 DGND 2.23e-19
C4427 DVDD.n47 DGND 9.76e-19
C4428 DVDD.t201 DGND 1.51e-19
C4429 DVDD.t493 DGND 1.51e-19
C4430 DVDD.n48 DGND 3.12e-19
C4431 DVDD.n49 DGND 0.001184f
C4432 DVDD.n50 DGND 0.00105f
C4433 DVDD.t348 DGND 0.001428f
C4434 DVDD.n51 DGND 0.001662f
C4435 DVDD.n52 DGND 0.001171f
C4436 DVDD.n53 DGND 4.15e-19
C4437 DVDD.n54 DGND 0.00105f
C4438 DVDD.n55 DGND 0.001892f
C4439 DVDD.t171 DGND 0.014144f
C4440 DVDD.t470 DGND 0.00605f
C4441 DVDD.t532 DGND 0.005794f
C4442 DVDD.t292 DGND 0.003579f
C4443 DVDD.t202 DGND 0.003579f
C4444 DVDD.t394 DGND 0.003579f
C4445 DVDD.t494 DGND 0.003579f
C4446 DVDD.t411 DGND 0.003579f
C4447 DVDD.t329 DGND 0.003579f
C4448 DVDD.t18 DGND 0.008009f
C4449 DVDD.t533 DGND 0.009628f
C4450 DVDD.t200 DGND 0.007157f
C4451 DVDD.t492 DGND 0.003962f
C4452 DVDD.t347 DGND 0.003792f
C4453 DVDD.t528 DGND 0.007498f
C4454 DVDD.t203 DGND 0.007157f
C4455 DVDD.t232 DGND 0.005411f
C4456 DVDD.n56 DGND 0.001231f
C4457 DVDD.t400 DGND 3.58e-19
C4458 DVDD.t250 DGND 3.58e-19
C4459 DVDD.n57 DGND 7.69e-19
C4460 DVDD.n58 DGND 8.77e-19
C4461 DVDD.n59 DGND 0.00105f
C4462 DVDD.t41 DGND 7.6e-19
C4463 DVDD.n60 DGND 4.15e-19
C4464 DVDD.n61 DGND 0.00105f
C4465 DVDD.t451 DGND 0.00156f
C4466 DVDD.n62 DGND 0.001598f
C4467 DVDD.n63 DGND 0.00105f
C4468 DVDD.t125 DGND 1.51e-19
C4469 DVDD.t256 DGND 1.51e-19
C4470 DVDD.n64 DGND 3.12e-19
C4471 DVDD.t164 DGND 5.49e-19
C4472 DVDD.n65 DGND 0.001052f
C4473 DVDD.n66 DGND 0.001415f
C4474 DVDD.t475 DGND 1.51e-19
C4475 DVDD.t179 DGND 1.51e-19
C4476 DVDD.n67 DGND 3.12e-19
C4477 DVDD.n68 DGND 4.15e-19
C4478 DVDD.n69 DGND 0.00105f
C4479 DVDD.t84 DGND 3.58e-19
C4480 DVDD.t154 DGND 3.58e-19
C4481 DVDD.n70 DGND 7.77e-19
C4482 DVDD.n71 DGND 3.75e-19
C4483 DVDD.n72 DGND 0.00105f
C4484 DVDD.t229 DGND 7.66e-19
C4485 DVDD.n73 DGND 0.001178f
C4486 DVDD.n74 DGND 0.001641f
C4487 DVDD.t345 DGND 7.6e-19
C4488 DVDD.n75 DGND 3.86e-19
C4489 DVDD.n76 DGND 0.001385f
C4490 DVDD.n77 DGND 0.002659f
C4491 DVDD.n78 DGND 0.003071f
C4492 DVDD.t518 DGND 0.001258f
C4493 DVDD.n79 DGND 7.9e-19
C4494 DVDD.n80 DGND 3.39e-19
C4495 DVDD.n81 DGND 0.00105f
C4496 DVDD.n82 DGND 0.00105f
C4497 DVDD.n83 DGND 2.62e-19
C4498 DVDD.n84 DGND 4.15e-19
C4499 DVDD.n85 DGND 0.00105f
C4500 DVDD.n86 DGND 0.00105f
C4501 DVDD.n87 DGND 0.00105f
C4502 DVDD.n88 DGND 2.12e-19
C4503 DVDD.n89 DGND 9.14e-19
C4504 DVDD.n90 DGND 4.99e-19
C4505 DVDD.n91 DGND 0.001377f
C4506 DVDD.n92 DGND 0.00105f
C4507 DVDD.n93 DGND 2.23e-19
C4508 DVDD.n94 DGND 9.76e-19
C4509 DVDD.n95 DGND 2.5e-19
C4510 DVDD.n96 DGND 2.32e-19
C4511 DVDD.n97 DGND 0.001552f
C4512 DVDD.n98 DGND 0.001377f
C4513 DVDD.t351 DGND 0.001428f
C4514 DVDD.n99 DGND 0.001171f
C4515 DVDD.n100 DGND 0.001662f
C4516 DVDD.n101 DGND 3.59e-19
C4517 DVDD.n102 DGND 0.00105f
C4518 DVDD.n103 DGND 0.00105f
C4519 DVDD.n104 DGND 2.3e-19
C4520 DVDD.n105 DGND 0.001184f
C4521 DVDD.n106 DGND 2.78e-19
C4522 DVDD.n107 DGND 4.15e-19
C4523 DVDD.n108 DGND 0.00137f
C4524 DVDD.n109 DGND 0.00105f
C4525 DVDD.n110 DGND 0.001517f
C4526 DVDD.n111 DGND 2.3e-19
C4527 DVDD.n112 DGND 3.45e-19
C4528 DVDD.n113 DGND 0.00105f
C4529 DVDD.n114 DGND 0.00105f
C4530 DVDD.n115 DGND 3.86e-19
C4531 DVDD.n116 DGND 0.001385f
C4532 DVDD.n117 DGND 0.00105f
C4533 DVDD.n118 DGND 0.00105f
C4534 DVDD.n119 DGND 3.41e-19
C4535 DVDD.t129 DGND 0.001429f
C4536 DVDD.n120 DGND 0.001838f
C4537 DVDD.n121 DGND 0.00263f
C4538 DVDD.n122 DGND 0.008232f
C4539 DVDD.t444 DGND 0.013548f
C4540 DVDD.n123 DGND 0.001253f
C4541 DVDD.t303 DGND 0.001428f
C4542 DVDD.n124 DGND 0.001662f
C4543 DVDD.n125 DGND 0.005448f
C4544 DVDD.n126 DGND 0.00137f
C4545 DVDD.n127 DGND 3.59e-19
C4546 DVDD.n128 DGND 0.001377f
C4547 DVDD.n129 DGND 0.001231f
C4548 DVDD.t445 DGND 0.001429f
C4549 DVDD.t305 DGND 3.58e-19
C4550 DVDD.t135 DGND 3.58e-19
C4551 DVDD.n130 DGND 7.69e-19
C4552 DVDD.n131 DGND 8.77e-19
C4553 DVDD.n132 DGND 0.00105f
C4554 DVDD.n133 DGND 4.15e-19
C4555 DVDD.n134 DGND 0.00105f
C4556 DVDD.n135 DGND 2.3e-19
C4557 DVDD.t320 DGND 0.00156f
C4558 DVDD.n136 DGND 0.001598f
C4559 DVDD.n137 DGND 2.3e-19
C4560 DVDD.n138 DGND 0.001171f
C4561 DVDD.n139 DGND 0.00105f
C4562 DVDD.t239 DGND 0.001428f
C4563 DVDD.n140 DGND 0.001662f
C4564 DVDD.n141 DGND 0.001415f
C4565 DVDD.t383 DGND 5.49e-19
C4566 DVDD.n142 DGND 0.001052f
C4567 DVDD.n143 DGND 4.15e-19
C4568 DVDD.n144 DGND 0.001377f
C4569 DVDD.n145 DGND 0.00105f
C4570 DVDD.t418 DGND 3.58e-19
C4571 DVDD.t425 DGND 3.58e-19
C4572 DVDD.n146 DGND 7.77e-19
C4573 DVDD.n147 DGND 3.75e-19
C4574 DVDD.n148 DGND 0.00105f
C4575 DVDD.t74 DGND 7.66e-19
C4576 DVDD.n149 DGND 0.001178f
C4577 DVDD.n150 DGND 0.001641f
C4578 DVDD.t362 DGND 0.001258f
C4579 DVDD.n151 DGND 7.9e-19
C4580 DVDD.n152 DGND 0.001892f
C4581 DVDD.n153 DGND 4.15e-19
C4582 DVDD.n154 DGND 0.001171f
C4583 DVDD.t107 DGND 1.51e-19
C4584 DVDD.t2 DGND 1.51e-19
C4585 DVDD.n155 DGND 3.12e-19
C4586 DVDD.n156 DGND 0.001184f
C4587 DVDD.n157 DGND 0.00105f
C4588 DVDD.t79 DGND 0.001428f
C4589 DVDD.n158 DGND 0.001662f
C4590 DVDD.n159 DGND 0.002427f
C4591 DVDD.t118 DGND 1.51e-19
C4592 DVDD.t459 DGND 1.51e-19
C4593 DVDD.n160 DGND 3.12e-19
C4594 DVDD.n161 DGND 9.76e-19
C4595 DVDD.n162 DGND 4.07e-19
C4596 DVDD.n163 DGND 2.23e-19
C4597 DVDD.n164 DGND 0.0021f
C4598 DVDD.t97 DGND 3.58e-19
C4599 DVDD.t288 DGND 3.58e-19
C4600 DVDD.n165 DGND 7.77e-19
C4601 DVDD.n166 DGND 0.001006f
C4602 DVDD.t368 DGND 0.001258f
C4603 DVDD.n167 DGND 4.12e-19
C4604 DVDD.n168 DGND 4.15e-19
C4605 DVDD.n169 DGND 4.15e-19
C4606 DVDD.n170 DGND 0.004927f
C4607 DVDD.n171 DGND 4.12e-19
C4608 DVDD.t64 DGND 7.66e-19
C4609 DVDD.n172 DGND 4.15e-19
C4610 DVDD.n173 DGND 0.0021f
C4611 DVDD.t387 DGND 0.001258f
C4612 DVDD.t116 DGND 3.58e-19
C4613 DVDD.t189 DGND 3.58e-19
C4614 DVDD.n174 DGND 7.77e-19
C4615 DVDD.n175 DGND 0.001006f
C4616 DVDD.n176 DGND 0.0021f
C4617 DVDD.t366 DGND 1.51e-19
C4618 DVDD.t103 DGND 1.51e-19
C4619 DVDD.n177 DGND 3.12e-19
C4620 DVDD.t416 DGND 5.49e-19
C4621 DVDD.n178 DGND 0.001052f
C4622 DVDD.n179 DGND 0.001377f
C4623 DVDD.n180 DGND 0.00105f
C4624 DVDD.t62 DGND 1.51e-19
C4625 DVDD.t212 DGND 1.51e-19
C4626 DVDD.n181 DGND 3.12e-19
C4627 DVDD.n182 DGND 4.15e-19
C4628 DVDD.n183 DGND 0.001253f
C4629 DVDD.t464 DGND 7.6e-19
C4630 DVDD.n184 DGND 0.001385f
C4631 DVDD.n185 DGND 0.002659f
C4632 DVDD.n186 DGND 0.00263f
C4633 DVDD.t407 DGND 0.014144f
C4634 DVDD.t138 DGND 0.00605f
C4635 DVDD.t335 DGND 0.005794f
C4636 DVDD.t306 DGND 0.003579f
C4637 DVDD.t272 DGND 0.003579f
C4638 DVDD.t27 DGND 0.003579f
C4639 DVDD.t515 DGND 0.003579f
C4640 DVDD.t166 DGND 0.003579f
C4641 DVDD.t502 DGND 0.003579f
C4642 DVDD.t93 DGND 0.008009f
C4643 DVDD.t14 DGND 0.009628f
C4644 DVDD.t270 DGND 0.007157f
C4645 DVDD.t140 DGND 0.003962f
C4646 DVDD.t195 DGND 0.003792f
C4647 DVDD.t241 DGND 0.007498f
C4648 DVDD.t269 DGND 0.007157f
C4649 DVDD.t246 DGND 0.005411f
C4650 DVDD.n187 DGND 0.001253f
C4651 DVDD.n188 DGND 0.00105f
C4652 DVDD.n189 DGND 3.39e-19
C4653 DVDD.n190 DGND 0.00105f
C4654 DVDD.n191 DGND 4.15e-19
C4655 DVDD.n192 DGND 0.00105f
C4656 DVDD.t523 DGND 0.001258f
C4657 DVDD.n193 DGND 7.9e-19
C4658 DVDD.t173 DGND 3.58e-19
C4659 DVDD.t343 DGND 3.58e-19
C4660 DVDD.n194 DGND 7.77e-19
C4661 DVDD.n195 DGND 9.14e-19
C4662 DVDD.n196 DGND 0.00105f
C4663 DVDD.t284 DGND 1.51e-19
C4664 DVDD.t454 DGND 1.51e-19
C4665 DVDD.n197 DGND 3.12e-19
C4666 DVDD.n198 DGND 9.76e-19
C4667 DVDD.n199 DGND 0.001552f
C4668 DVDD.t486 DGND 1.51e-19
C4669 DVDD.t276 DGND 1.51e-19
C4670 DVDD.n200 DGND 3.12e-19
C4671 DVDD.n201 DGND 0.001184f
C4672 DVDD.n202 DGND 0.001377f
C4673 DVDD.n203 DGND 0.00105f
C4674 DVDD.t322 DGND 0.001428f
C4675 DVDD.n204 DGND 0.00137f
C4676 DVDD.n205 DGND 3.86e-19
C4677 DVDD.n206 DGND 0.00105f
C4678 DVDD.n207 DGND 0.00105f
C4679 DVDD.t199 DGND 0.00156f
C4680 DVDD.n208 DGND 0.001517f
C4681 DVDD.t527 DGND 3.58e-19
C4682 DVDD.t224 DGND 3.58e-19
C4683 DVDD.n209 DGND 7.69e-19
C4684 DVDD.n210 DGND 8.77e-19
C4685 DVDD.t509 DGND 0.001429f
C4686 DVDD.n211 DGND 0.001838f
C4687 DVDD.n212 DGND 3.41e-19
C4688 DVDD.n213 DGND 0.00105f
C4689 DVDD.n214 DGND 0.001231f
C4690 DVDD.t286 DGND 7.6e-19
C4691 DVDD.n215 DGND 0.001385f
C4692 DVDD.n216 DGND 0.00105f
C4693 DVDD.n217 DGND 0.00105f
C4694 DVDD.n218 DGND 2.3e-19
C4695 DVDD.n219 DGND 3.45e-19
C4696 DVDD.n220 DGND 0.00105f
C4697 DVDD.n221 DGND 0.00105f
C4698 DVDD.n222 DGND 4.15e-19
C4699 DVDD.n223 DGND 4.15e-19
C4700 DVDD.n224 DGND 2.78e-19
C4701 DVDD.n225 DGND 0.001598f
C4702 DVDD.n226 DGND 0.001171f
C4703 DVDD.n227 DGND 0.001662f
C4704 DVDD.n228 DGND 3.59e-19
C4705 DVDD.n229 DGND 0.00105f
C4706 DVDD.n230 DGND 0.00105f
C4707 DVDD.n231 DGND 2.3e-19
C4708 DVDD.t439 DGND 5.49e-19
C4709 DVDD.n232 DGND 0.001052f
C4710 DVDD.n233 DGND 2.32e-19
C4711 DVDD.n234 DGND 2.5e-19
C4712 DVDD.n235 DGND 0.001415f
C4713 DVDD.n236 DGND 4.99e-19
C4714 DVDD.n237 DGND 0.001377f
C4715 DVDD.n238 DGND 0.00105f
C4716 DVDD.n239 DGND 2.23e-19
C4717 DVDD.n240 DGND 4.15e-19
C4718 DVDD.n241 DGND 0.00105f
C4719 DVDD.n242 DGND 0.00105f
C4720 DVDD.n243 DGND 2.12e-19
C4721 DVDD.n244 DGND 3.75e-19
C4722 DVDD.n245 DGND 0.00105f
C4723 DVDD.n246 DGND 0.00105f
C4724 DVDD.n247 DGND 2.62e-19
C4725 DVDD.t278 DGND 7.66e-19
C4726 DVDD.n248 DGND 0.001178f
C4727 DVDD.n249 DGND 0.001641f
C4728 DVDD.n250 DGND 0.003071f
C4729 DVDD.t99 DGND 7.6e-19
C4730 DVDD.n251 DGND 4.15e-19
C4731 DVDD.n252 DGND 0.00105f
C4732 DVDD.n253 DGND 0.001377f
C4733 DVDD.n254 DGND 2.78e-19
C4734 DVDD.t271 DGND 1.51e-19
C4735 DVDD.t141 DGND 1.51e-19
C4736 DVDD.n255 DGND 3.12e-19
C4737 DVDD.t15 DGND 5.49e-19
C4738 DVDD.n256 DGND 0.001052f
C4739 DVDD.n257 DGND 2.32e-19
C4740 DVDD.t28 DGND 3.58e-19
C4741 DVDD.t167 DGND 3.58e-19
C4742 DVDD.n258 DGND 7.77e-19
C4743 DVDD.n259 DGND 0.001006f
C4744 DVDD.n260 DGND 0.0021f
C4745 DVDD.t516 DGND 1.51e-19
C4746 DVDD.t503 DGND 1.51e-19
C4747 DVDD.n261 DGND 3.12e-19
C4748 DVDD.n262 DGND 4.15e-19
C4749 DVDD.n263 DGND 0.0021f
C4750 DVDD.t307 DGND 0.001258f
C4751 DVDD.t82 DGND 0.001258f
C4752 DVDD.n264 DGND 9.69e-19
C4753 DVDD.n265 DGND 0.00135f
C4754 DVDD.t45 DGND 3.58e-19
C4755 DVDD.t274 DGND 3.58e-19
C4756 DVDD.n266 DGND 7.77e-19
C4757 DVDD.n267 DGND 0.003693f
C4758 DVDD.t257 DGND 0.009969f
C4759 DVDD.t81 DGND 0.005794f
C4760 DVDD.t44 DGND 0.003579f
C4761 DVDD.t273 DGND 0.003579f
C4762 DVDD.t67 DGND 0.008584f
C4763 DVDD.t242 DGND 0.013249f
C4764 DVDD.t491 DGND 0.009969f
C4765 DVDD.t481 DGND 0.005794f
C4766 DVDD.t100 DGND 0.003579f
C4767 DVDD.t121 DGND 0.003579f
C4768 DVDD.t519 DGND 0.008584f
C4769 DVDD.t24 DGND 0.013249f
C4770 DVDD.t59 DGND 0.001258f
C4771 DVDD.n268 DGND 9.69e-19
C4772 DVDD.n269 DGND 0.00135f
C4773 DVDD.t88 DGND 3.58e-19
C4774 DVDD.t92 DGND 3.58e-19
C4775 DVDD.n270 DGND 7.77e-19
C4776 DVDD.t5 DGND 2.06e-19
C4777 DVDD.t147 DGND 1.62e-19
C4778 DVDD.n271 DGND 3.98e-19
C4779 DVDD.n272 DGND 9.86e-19
C4780 DVDD.n273 DGND 0.001172f
C4781 DVDD.n274 DGND 4.15e-19
C4782 DVDD.n275 DGND 0.001172f
C4783 DVDD.t149 DGND 2.94e-19
C4784 DVDD.t52 DGND 9.54e-20
C4785 DVDD.n276 DGND 0.001417f
C4786 DVDD.n277 DGND 0.001172f
C4787 DVDD.t191 DGND 2.94e-19
C4788 DVDD.t327 DGND 9.54e-20
C4789 DVDD.n278 DGND 0.001417f
C4790 DVDD.n279 DGND 4.15e-19
C4791 DVDD.n280 DGND 0.001172f
C4792 DVDD.t193 DGND 1.62e-19
C4793 DVDD.t231 DGND 2.06e-19
C4794 DVDD.n281 DGND 3.98e-19
C4795 DVDD.n282 DGND 9.86e-19
C4796 DVDD.t282 DGND 3.58e-19
C4797 DVDD.t280 DGND 3.58e-19
C4798 DVDD.n283 DGND 7.77e-19
C4799 DVDD.n284 DGND 0.001006f
C4800 DVDD.n285 DGND 0.001412f
C4801 DVDD.t299 DGND 0.001258f
C4802 DVDD.n286 DGND 9.69e-19
C4803 DVDD.n287 DGND 3.75e-19
C4804 DVDD.n288 DGND 2.12e-19
C4805 DVDD.n289 DGND 0.00135f
C4806 DVDD.n290 DGND 0.003854f
C4807 DVDD.t264 DGND 0.001489f
C4808 DVDD.n291 DGND 0.00658f
C4809 DVDD.n292 DGND 0.003099f
C4810 DVDD.n293 DGND 0.00135f
C4811 DVDD.n294 DGND 3.11e-19
C4812 DVDD.n295 DGND 4.15e-19
C4813 DVDD.n296 DGND 4.15e-19
C4814 DVDD.n297 DGND 0.001172f
C4815 DVDD.n298 DGND 0.001172f
C4816 DVDD.n299 DGND 0.001172f
C4817 DVDD.n300 DGND 4.15e-19
C4818 DVDD.n301 DGND 2.12e-19
C4819 DVDD.n302 DGND 0.0012f
C4820 DVDD.n303 DGND 0.001979f
C4821 DVDD.n304 DGND 0.001979f
C4822 DVDD.n305 DGND 0.0012f
C4823 DVDD.n306 DGND 2.12e-19
C4824 DVDD.n307 DGND 4.15e-19
C4825 DVDD.n308 DGND 0.001172f
C4826 DVDD.n309 DGND 0.001172f
C4827 DVDD.n310 DGND 0.001172f
C4828 DVDD.n311 DGND 4.15e-19
C4829 DVDD.n312 DGND 4.15e-19
C4830 DVDD.n313 DGND 3.11e-19
C4831 DVDD.n314 DGND 0.00135f
C4832 DVDD.n315 DGND 0.003099f
C4833 DVDD.t462 DGND 0.001489f
C4834 DVDD.n316 DGND 0.00658f
C4835 DVDD.n317 DGND 0.003854f
C4836 DVDD.n318 DGND 0.001006f
C4837 DVDD.n319 DGND 2.12e-19
C4838 DVDD.n320 DGND 3.75e-19
C4839 DVDD.n321 DGND 0.001412f
C4840 DVDD.n322 DGND 0.003693f
C4841 DVDD.t122 DGND 3.58e-19
C4842 DVDD.t101 DGND 3.58e-19
C4843 DVDD.n323 DGND 7.77e-19
C4844 DVDD.n324 DGND 0.001006f
C4845 DVDD.n325 DGND 0.001412f
C4846 DVDD.t482 DGND 0.001258f
C4847 DVDD.n326 DGND 9.69e-19
C4848 DVDD.n327 DGND 3.75e-19
C4849 DVDD.n328 DGND 2.12e-19
C4850 DVDD.n329 DGND 0.00135f
C4851 DVDD.n330 DGND 0.003854f
C4852 DVDD.t25 DGND 0.001489f
C4853 DVDD.n331 DGND 0.006355f
C4854 DVDD.n332 DGND 0.006566f
C4855 DVDD.n333 DGND 0.013469f
C4856 DVDD.t376 DGND 0.009756f
C4857 DVDD.t58 DGND 0.005794f
C4858 DVDD.t91 DGND 0.003579f
C4859 DVDD.t87 DGND 0.003579f
C4860 DVDD.t60 DGND 0.008584f
C4861 DVDD.t461 DGND 0.014272f
C4862 DVDD.t146 DGND 0.009522f
C4863 DVDD.t4 DGND 0.003579f
C4864 DVDD.t457 DGND 0.006092f
C4865 DVDD.t220 DGND 0.006752f
C4866 DVDD.t148 DGND 0.004516f
C4867 DVDD.t51 DGND 0.007945f
C4868 DVDD.t326 DGND 0.007945f
C4869 DVDD.t190 DGND 0.004516f
C4870 DVDD.t46 DGND 0.006752f
C4871 DVDD.t162 DGND 0.006092f
C4872 DVDD.t230 DGND 0.003579f
C4873 DVDD.t192 DGND 0.009522f
C4874 DVDD.t263 DGND 0.014272f
C4875 DVDD.t7 DGND 0.008584f
C4876 DVDD.t279 DGND 0.003579f
C4877 DVDD.t281 DGND 0.003579f
C4878 DVDD.t298 DGND 0.005794f
C4879 DVDD.t358 DGND 0.009756f
C4880 DVDD.n334 DGND 0.013469f
C4881 DVDD.n335 DGND 0.006566f
C4882 DVDD.t243 DGND 0.001489f
C4883 DVDD.n336 DGND 0.006355f
C4884 DVDD.n337 DGND 0.003854f
C4885 DVDD.n338 DGND 0.001006f
C4886 DVDD.n339 DGND 2.12e-19
C4887 DVDD.n340 DGND 3.75e-19
C4888 DVDD.n341 DGND 0.001412f
C4889 DVDD.n342 DGND 0.004927f
C4890 DVDD.n343 DGND 0.018475f
C4891 DVDD.n344 DGND 0.002811f
C4892 DVDD.t139 DGND 7.66e-19
C4893 DVDD.n345 DGND 0.001178f
C4894 DVDD.n346 DGND 2.62e-19
C4895 DVDD.n347 DGND 0.0021f
C4896 DVDD.n348 DGND 4.12e-19
C4897 DVDD.n349 DGND 3.39e-19
C4898 DVDD.n350 DGND 7.9e-19
C4899 DVDD.n351 DGND 2.12e-19
C4900 DVDD.n352 DGND 3.75e-19
C4901 DVDD.n353 DGND 0.0021f
C4902 DVDD.n354 DGND 4.15e-19
C4903 DVDD.n355 DGND 2.23e-19
C4904 DVDD.n356 DGND 9.76e-19
C4905 DVDD.n357 DGND 2.5e-19
C4906 DVDD.n358 DGND 0.0021f
C4907 DVDD.n359 DGND 4.07e-19
C4908 DVDD.n360 DGND 0.002427f
C4909 DVDD.n361 DGND 0.001918f
C4910 DVDD.n362 DGND 2.3e-19
C4911 DVDD.n363 DGND 0.001184f
C4912 DVDD.n364 DGND 0.00105f
C4913 DVDD.n365 DGND 0.00105f
C4914 DVDD.n366 DGND 3.59e-19
C4915 DVDD.t196 DGND 0.001428f
C4916 DVDD.n367 DGND 0.001662f
C4917 DVDD.n368 DGND 0.001171f
C4918 DVDD.n369 DGND 0.001233f
C4919 DVDD.n370 DGND 0.001735f
C4920 DVDD.n371 DGND 4.15e-19
C4921 DVDD.n372 DGND 3.86e-19
C4922 DVDD.n373 DGND 0.001385f
C4923 DVDD.n374 DGND 0.002659f
C4924 DVDD.n375 DGND 0.001892f
C4925 DVDD.n376 DGND 0.001919f
C4926 DVDD.n377 DGND 0.005247f
C4927 DVDD.t98 DGND 0.011503f
C4928 DVDD.t490 DGND 0.017254f
C4929 DVDD.t277 DGND 0.008009f
C4930 DVDD.t522 DGND 0.003834f
C4931 DVDD.t452 DGND 0.003579f
C4932 DVDD.t172 DGND 0.003579f
C4933 DVDD.t487 DGND 0.003579f
C4934 DVDD.t342 DGND 0.003579f
C4935 DVDD.t283 DGND 0.003579f
C4936 DVDD.t514 DGND 0.003579f
C4937 DVDD.t453 DGND 0.011332f
C4938 DVDD.t438 DGND 0.010267f
C4939 DVDD.t321 DGND 0.003579f
C4940 DVDD.t485 DGND 0.004899f
C4941 DVDD.t275 DGND 0.00737f
C4942 DVDD.t262 DGND 0.007882f
C4943 DVDD.t484 DGND 0.004644f
C4944 DVDD.t198 DGND 0.003067f
C4945 DVDD.t37 DGND 0.00409f
C4946 DVDD.t526 DGND 0.00409f
C4947 DVDD.t285 DGND 0.003579f
C4948 DVDD.t223 DGND 0.004644f
C4949 DVDD.t508 DGND 0.017855f
C4950 DVDD.n378 DGND 0.018343f
C4951 DVDD.n379 DGND 0.001231f
C4952 DVDD.t301 DGND 0.001429f
C4953 DVDD.t456 DGND 3.58e-19
C4954 DVDD.t507 DGND 3.58e-19
C4955 DVDD.n380 DGND 7.69e-19
C4956 DVDD.n381 DGND 8.77e-19
C4957 DVDD.n382 DGND 0.00105f
C4958 DVDD.n383 DGND 4.15e-19
C4959 DVDD.n384 DGND 0.00105f
C4960 DVDD.n385 DGND 2.3e-19
C4961 DVDD.t469 DGND 0.00156f
C4962 DVDD.n386 DGND 0.001598f
C4963 DVDD.n387 DGND 2.3e-19
C4964 DVDD.n388 DGND 0.001171f
C4965 DVDD.n389 DGND 0.00105f
C4966 DVDD.t216 DGND 0.001428f
C4967 DVDD.n390 DGND 0.001662f
C4968 DVDD.n391 DGND 0.001415f
C4969 DVDD.t414 DGND 5.49e-19
C4970 DVDD.n392 DGND 0.001052f
C4971 DVDD.n393 DGND 4.15e-19
C4972 DVDD.n394 DGND 0.001377f
C4973 DVDD.n395 DGND 0.00105f
C4974 DVDD.t372 DGND 3.58e-19
C4975 DVDD.t32 DGND 3.58e-19
C4976 DVDD.n396 DGND 7.77e-19
C4977 DVDD.n397 DGND 3.75e-19
C4978 DVDD.n398 DGND 0.00105f
C4979 DVDD.t389 DGND 7.66e-19
C4980 DVDD.n399 DGND 0.001178f
C4981 DVDD.n400 DGND 0.001641f
C4982 DVDD.t385 DGND 0.001258f
C4983 DVDD.n401 DGND 7.9e-19
C4984 DVDD.n402 DGND 0.003071f
C4985 DVDD.n403 DGND 3.39e-19
C4986 DVDD.n404 DGND 0.00105f
C4987 DVDD.n405 DGND 0.00105f
C4988 DVDD.n406 DGND 2.62e-19
C4989 DVDD.n407 DGND 4.15e-19
C4990 DVDD.n408 DGND 0.00105f
C4991 DVDD.n409 DGND 0.00105f
C4992 DVDD.n410 DGND 2.12e-19
C4993 DVDD.n411 DGND 9.14e-19
C4994 DVDD.n412 DGND 4.99e-19
C4995 DVDD.n413 DGND 0.00105f
C4996 DVDD.n414 DGND 0.00105f
C4997 DVDD.n415 DGND 2.23e-19
C4998 DVDD.t339 DGND 1.51e-19
C4999 DVDD.t441 DGND 1.51e-19
C5000 DVDD.n416 DGND 3.12e-19
C5001 DVDD.n417 DGND 9.76e-19
C5002 DVDD.n418 DGND 2.5e-19
C5003 DVDD.n419 DGND 2.32e-19
C5004 DVDD.n420 DGND 0.001552f
C5005 DVDD.n421 DGND 0.001377f
C5006 DVDD.n422 DGND 3.59e-19
C5007 DVDD.n423 DGND 0.00105f
C5008 DVDD.n424 DGND 0.00105f
C5009 DVDD.t443 DGND 1.51e-19
C5010 DVDD.t21 DGND 1.51e-19
C5011 DVDD.n425 DGND 3.12e-19
C5012 DVDD.n426 DGND 0.001184f
C5013 DVDD.n427 DGND 2.78e-19
C5014 DVDD.n428 DGND 4.15e-19
C5015 DVDD.n429 DGND 0.00137f
C5016 DVDD.n430 DGND 0.00105f
C5017 DVDD.n431 DGND 0.001517f
C5018 DVDD.n432 DGND 3.45e-19
C5019 DVDD.n433 DGND 0.00105f
C5020 DVDD.n434 DGND 0.00105f
C5021 DVDD.n435 DGND 3.86e-19
C5022 DVDD.t90 DGND 7.6e-19
C5023 DVDD.n436 DGND 0.001385f
C5024 DVDD.n437 DGND 0.00105f
C5025 DVDD.n438 DGND 0.00105f
C5026 DVDD.n439 DGND 3.41e-19
C5027 DVDD.n440 DGND 0.001838f
C5028 DVDD.n441 DGND 0.00263f
C5029 DVDD.n442 DGND 0.018343f
C5030 DVDD.t300 DGND 0.017855f
C5031 DVDD.t455 DGND 0.004644f
C5032 DVDD.t89 DGND 0.003579f
C5033 DVDD.t506 DGND 0.00409f
C5034 DVDD.t197 DGND 0.00409f
C5035 DVDD.t468 DGND 0.003067f
C5036 DVDD.t22 DGND 0.004644f
C5037 DVDD.t460 DGND 0.007882f
C5038 DVDD.t442 DGND 0.00737f
C5039 DVDD.t20 DGND 0.004899f
C5040 DVDD.t215 DGND 0.003579f
C5041 DVDD.t413 DGND 0.010267f
C5042 DVDD.t338 DGND 0.011332f
C5043 DVDD.t289 DGND 0.003579f
C5044 DVDD.t440 DGND 0.003579f
C5045 DVDD.t371 DGND 0.003579f
C5046 DVDD.t23 DGND 0.003579f
C5047 DVDD.t31 DGND 0.003579f
C5048 DVDD.t401 DGND 0.003579f
C5049 DVDD.t384 DGND 0.003834f
C5050 DVDD.t388 DGND 0.008009f
C5051 DVDD.t222 DGND 0.017254f
C5052 DVDD.t463 DGND 0.011503f
C5053 DVDD.t313 DGND 0.014144f
C5054 DVDD.t63 DGND 0.00605f
C5055 DVDD.t13 DGND 0.005794f
C5056 DVDD.t386 DGND 0.003579f
C5057 DVDD.t210 DGND 0.003579f
C5058 DVDD.t188 DGND 0.003579f
C5059 DVDD.t102 DGND 0.003579f
C5060 DVDD.t115 DGND 0.003579f
C5061 DVDD.t365 DGND 0.003579f
C5062 DVDD.t159 DGND 0.008009f
C5063 DVDD.t415 DGND 0.009628f
C5064 DVDD.t211 DGND 0.007157f
C5065 DVDD.t61 DGND 0.003962f
C5066 DVDD.t314 DGND 0.003792f
C5067 DVDD.t26 DGND 0.007498f
C5068 DVDD.t213 DGND 0.007157f
C5069 DVDD.t483 DGND 0.005411f
C5070 DVDD.n443 DGND 0.005247f
C5071 DVDD.n444 DGND 0.001919f
C5072 DVDD.n445 DGND 0.001892f
C5073 DVDD.n446 DGND 0.00105f
C5074 DVDD.n447 DGND 3.86e-19
C5075 DVDD.n448 DGND 4.15e-19
C5076 DVDD.n449 DGND 0.001735f
C5077 DVDD.n450 DGND 0.001233f
C5078 DVDD.n451 DGND 0.001171f
C5079 DVDD.t315 DGND 0.001428f
C5080 DVDD.n452 DGND 0.001662f
C5081 DVDD.n453 DGND 3.59e-19
C5082 DVDD.n454 DGND 0.00105f
C5083 DVDD.n455 DGND 0.00105f
C5084 DVDD.n456 DGND 2.78e-19
C5085 DVDD.n457 DGND 0.001184f
C5086 DVDD.n458 DGND 2.3e-19
C5087 DVDD.n459 DGND 0.001918f
C5088 DVDD.n460 DGND 4.07e-19
C5089 DVDD.n461 DGND 0.002427f
C5090 DVDD.n462 DGND 2.32e-19
C5091 DVDD.n463 DGND 2.5e-19
C5092 DVDD.n464 DGND 9.76e-19
C5093 DVDD.n465 DGND 4.15e-19
C5094 DVDD.n466 DGND 2.23e-19
C5095 DVDD.n467 DGND 0.0021f
C5096 DVDD.n468 DGND 2.12e-19
C5097 DVDD.n469 DGND 3.75e-19
C5098 DVDD.n470 DGND 7.9e-19
C5099 DVDD.n471 DGND 3.39e-19
C5100 DVDD.n472 DGND 0.0021f
C5101 DVDD.n473 DGND 0.0021f
C5102 DVDD.n474 DGND 2.62e-19
C5103 DVDD.n475 DGND 0.001178f
C5104 DVDD.n476 DGND 0.002811f
C5105 DVDD.n477 DGND 0.018475f
C5106 DVDD.n478 DGND 4.12e-19
C5107 DVDD.t521 DGND 7.66e-19
C5108 DVDD.n479 DGND 4.15e-19
C5109 DVDD.n480 DGND 0.0021f
C5110 DVDD.t409 DGND 0.001258f
C5111 DVDD.t185 DGND 3.58e-19
C5112 DVDD.t109 DGND 3.58e-19
C5113 DVDD.n481 DGND 7.77e-19
C5114 DVDD.n482 DGND 0.001006f
C5115 DVDD.n483 DGND 0.0021f
C5116 DVDD.t183 DGND 1.51e-19
C5117 DVDD.t466 DGND 1.51e-19
C5118 DVDD.n484 DGND 3.12e-19
C5119 DVDD.t158 DGND 5.49e-19
C5120 DVDD.n485 DGND 0.001052f
C5121 DVDD.n486 DGND 0.001377f
C5122 DVDD.n487 DGND 0.00105f
C5123 DVDD.t500 DGND 1.51e-19
C5124 DVDD.t219 DGND 1.51e-19
C5125 DVDD.n488 DGND 3.12e-19
C5126 DVDD.n489 DGND 4.15e-19
C5127 DVDD.n490 DGND 0.001253f
C5128 DVDD.t437 DGND 7.6e-19
C5129 DVDD.n491 DGND 0.001385f
C5130 DVDD.n492 DGND 0.002659f
C5131 DVDD.t356 DGND 0.005656f
C5132 DVDD.n493 DGND 0.001253f
C5133 DVDD.n494 DGND 0.00105f
C5134 DVDD.n495 DGND 0.00137f
C5135 DVDD.t357 DGND 2.94e-19
C5136 DVDD.t120 DGND 9.54e-20
C5137 DVDD.n496 DGND 0.001417f
C5138 DVDD.n497 DGND 0.0012f
C5139 DVDD.n498 DGND 0.001552f
C5140 DVDD.t447 DGND 2.94e-19
C5141 DVDD.t378 DGND 9.54e-20
C5142 DVDD.n499 DGND 0.001417f
C5143 DVDD.n500 DGND 4.15e-19
C5144 DVDD.n501 DGND 0.001253f
C5145 DVDD.t170 DGND 0.014144f
C5146 DVDD.t29 DGND 0.00605f
C5147 DVDD.t312 DGND 0.005794f
C5148 DVDD.t488 DGND 0.003579f
C5149 DVDD.t50 DGND 0.003579f
C5150 DVDD.t472 DGND 0.003579f
C5151 DVDD.t168 DGND 0.003579f
C5152 DVDD.t391 DGND 0.003579f
C5153 DVDD.t233 DGND 0.003579f
C5154 DVDD.t53 DGND 0.008009f
C5155 DVDD.t235 DGND 0.009628f
C5156 DVDD.t48 DGND 0.007157f
C5157 DVDD.t10 DGND 0.003962f
C5158 DVDD.t529 DGND 0.003792f
C5159 DVDD.t194 DGND 0.007498f
C5160 DVDD.t47 DGND 0.007157f
C5161 DVDD.t72 DGND 0.005411f
C5162 DVDD.n502 DGND 0.001253f
C5163 DVDD.n503 DGND 0.00105f
C5164 DVDD.n504 DGND 3.39e-19
C5165 DVDD.n505 DGND 0.00105f
C5166 DVDD.n506 DGND 4.15e-19
C5167 DVDD.n507 DGND 0.00105f
C5168 DVDD.t77 DGND 0.001258f
C5169 DVDD.n508 DGND 7.9e-19
C5170 DVDD.t341 DGND 3.58e-19
C5171 DVDD.t227 DGND 3.58e-19
C5172 DVDD.n509 DGND 7.77e-19
C5173 DVDD.n510 DGND 9.14e-19
C5174 DVDD.n511 DGND 0.00105f
C5175 DVDD.t57 DGND 1.51e-19
C5176 DVDD.t525 DGND 1.51e-19
C5177 DVDD.n512 DGND 3.12e-19
C5178 DVDD.n513 DGND 9.76e-19
C5179 DVDD.n514 DGND 0.001552f
C5180 DVDD.t260 DGND 1.51e-19
C5181 DVDD.t332 DGND 1.51e-19
C5182 DVDD.n515 DGND 3.12e-19
C5183 DVDD.n516 DGND 0.001184f
C5184 DVDD.n517 DGND 0.001377f
C5185 DVDD.n518 DGND 0.00105f
C5186 DVDD.t112 DGND 0.001428f
C5187 DVDD.n519 DGND 0.00137f
C5188 DVDD.n520 DGND 3.86e-19
C5189 DVDD.n521 DGND 0.001377f
C5190 DVDD.n522 DGND 0.00105f
C5191 DVDD.t449 DGND 1.62e-19
C5192 DVDD.t511 DGND 2.06e-19
C5193 DVDD.n523 DGND 3.98e-19
C5194 DVDD.n524 DGND 4.15e-19
C5195 DVDD.n525 DGND 0.00105f
C5196 DVDD.n526 DGND 0.001598f
C5197 DVDD.n527 DGND 4.15e-19
C5198 DVDD.n528 DGND 0.00137f
C5199 DVDD.n529 DGND 0.001231f
C5200 DVDD.t360 DGND 7.6e-19
C5201 DVDD.n530 DGND 0.001385f
C5202 DVDD.n531 DGND 0.00105f
C5203 DVDD.n532 DGND 0.00105f
C5204 DVDD.n533 DGND 3.11e-19
C5205 DVDD.n534 DGND 8.64e-19
C5206 DVDD.n535 DGND 3.99e-19
C5207 DVDD.n536 DGND 0.00105f
C5208 DVDD.n537 DGND 0.00105f
C5209 DVDD.n538 DGND 4.15e-19
C5210 DVDD.n539 DGND 4.15e-19
C5211 DVDD.n540 DGND 2.78e-19
C5212 DVDD.n541 DGND 0.001598f
C5213 DVDD.n542 DGND 0.001171f
C5214 DVDD.n543 DGND 0.001662f
C5215 DVDD.n544 DGND 3.59e-19
C5216 DVDD.n545 DGND 0.00105f
C5217 DVDD.n546 DGND 0.00105f
C5218 DVDD.n547 DGND 2.3e-19
C5219 DVDD.t513 DGND 5.49e-19
C5220 DVDD.n548 DGND 0.001052f
C5221 DVDD.n549 DGND 2.32e-19
C5222 DVDD.n550 DGND 2.5e-19
C5223 DVDD.n551 DGND 0.001415f
C5224 DVDD.n552 DGND 4.99e-19
C5225 DVDD.n553 DGND 0.001377f
C5226 DVDD.n554 DGND 0.00105f
C5227 DVDD.n555 DGND 2.23e-19
C5228 DVDD.n556 DGND 4.15e-19
C5229 DVDD.n557 DGND 0.00105f
C5230 DVDD.n558 DGND 0.00105f
C5231 DVDD.n559 DGND 2.12e-19
C5232 DVDD.n560 DGND 3.75e-19
C5233 DVDD.n561 DGND 0.00105f
C5234 DVDD.n562 DGND 0.00105f
C5235 DVDD.n563 DGND 2.62e-19
C5236 DVDD.t403 DGND 7.66e-19
C5237 DVDD.n564 DGND 0.001178f
C5238 DVDD.n565 DGND 0.001641f
C5239 DVDD.n566 DGND 0.003071f
C5240 DVDD.t66 DGND 7.6e-19
C5241 DVDD.n567 DGND 4.15e-19
C5242 DVDD.n568 DGND 0.00105f
C5243 DVDD.n569 DGND 0.001377f
C5244 DVDD.n570 DGND 2.78e-19
C5245 DVDD.t49 DGND 1.51e-19
C5246 DVDD.t11 DGND 1.51e-19
C5247 DVDD.n571 DGND 3.12e-19
C5248 DVDD.t236 DGND 5.49e-19
C5249 DVDD.n572 DGND 0.001052f
C5250 DVDD.n573 DGND 2.32e-19
C5251 DVDD.t473 DGND 3.58e-19
C5252 DVDD.t392 DGND 3.58e-19
C5253 DVDD.n574 DGND 7.77e-19
C5254 DVDD.n575 DGND 0.001006f
C5255 DVDD.n576 DGND 0.0021f
C5256 DVDD.t169 DGND 1.51e-19
C5257 DVDD.t234 DGND 1.51e-19
C5258 DVDD.n577 DGND 3.12e-19
C5259 DVDD.n578 DGND 4.15e-19
C5260 DVDD.n579 DGND 0.0021f
C5261 DVDD.t489 DGND 0.001258f
C5262 DVDD.n580 DGND 0.002811f
C5263 DVDD.t30 DGND 7.66e-19
C5264 DVDD.n581 DGND 0.001178f
C5265 DVDD.n582 DGND 2.62e-19
C5266 DVDD.n583 DGND 0.0021f
C5267 DVDD.n584 DGND 4.12e-19
C5268 DVDD.n585 DGND 3.39e-19
C5269 DVDD.n586 DGND 7.9e-19
C5270 DVDD.n587 DGND 2.12e-19
C5271 DVDD.n588 DGND 3.75e-19
C5272 DVDD.n589 DGND 0.0021f
C5273 DVDD.n590 DGND 4.15e-19
C5274 DVDD.n591 DGND 2.23e-19
C5275 DVDD.n592 DGND 9.76e-19
C5276 DVDD.n593 DGND 2.5e-19
C5277 DVDD.n594 DGND 0.0021f
C5278 DVDD.n595 DGND 4.07e-19
C5279 DVDD.n596 DGND 0.002427f
C5280 DVDD.n597 DGND 0.001918f
C5281 DVDD.n598 DGND 2.3e-19
C5282 DVDD.n599 DGND 0.001184f
C5283 DVDD.n600 DGND 0.00105f
C5284 DVDD.n601 DGND 0.00105f
C5285 DVDD.n602 DGND 3.59e-19
C5286 DVDD.t530 DGND 0.001428f
C5287 DVDD.n603 DGND 0.001662f
C5288 DVDD.n604 DGND 0.001171f
C5289 DVDD.n605 DGND 0.001233f
C5290 DVDD.n606 DGND 0.001735f
C5291 DVDD.n607 DGND 4.15e-19
C5292 DVDD.n608 DGND 3.86e-19
C5293 DVDD.n609 DGND 0.001385f
C5294 DVDD.n610 DGND 0.002659f
C5295 DVDD.n611 DGND 0.001892f
C5296 DVDD.n612 DGND 0.001919f
C5297 DVDD.n613 DGND 0.005247f
C5298 DVDD.t65 DGND 0.011503f
C5299 DVDD.t136 DGND 0.017254f
C5300 DVDD.t402 DGND 0.008009f
C5301 DVDD.t76 DGND 0.003834f
C5302 DVDD.t290 DGND 0.003579f
C5303 DVDD.t340 DGND 0.003579f
C5304 DVDD.t261 DGND 0.003579f
C5305 DVDD.t226 DGND 0.003579f
C5306 DVDD.t56 DGND 0.003579f
C5307 DVDD.t237 DGND 0.003579f
C5308 DVDD.t524 DGND 0.011332f
C5309 DVDD.t512 DGND 0.010267f
C5310 DVDD.t111 DGND 0.003579f
C5311 DVDD.t259 DGND 0.004899f
C5312 DVDD.t331 DGND 0.00737f
C5313 DVDD.t323 DGND 0.007882f
C5314 DVDD.t258 DGND 0.006263f
C5315 DVDD.t448 DGND 0.003067f
C5316 DVDD.t328 DGND 0.00409f
C5317 DVDD.t510 DGND 0.00409f
C5318 DVDD.t359 DGND 0.003067f
C5319 DVDD.t297 DGND 0.01129f
C5320 DVDD.t479 DGND 0.01244f
C5321 DVDD.t119 DGND 0.01015f
C5322 DVDD.t377 DGND 0.01015f
C5323 DVDD.t446 DGND 0.005656f
C5324 DVDD.n614 DGND 0.005545f
C5325 DVDD.n615 DGND 0.001919f
C5326 DVDD.n616 DGND 0.001253f
C5327 DVDD.n617 DGND 0.00105f
C5328 DVDD.n618 DGND 4.15e-19
C5329 DVDD.n619 DGND 2.12e-19
C5330 DVDD.n620 DGND 0.0012f
C5331 DVDD.n621 DGND 0.00329f
C5332 DVDD.n622 DGND 0.00329f
C5333 DVDD.n623 DGND 0.001552f
C5334 DVDD.n624 DGND 2.12e-19
C5335 DVDD.n625 DGND 4.15e-19
C5336 DVDD.n626 DGND 3.11e-19
C5337 DVDD.n627 DGND 0.001231f
C5338 DVDD.n628 DGND 0.00105f
C5339 DVDD.n629 DGND 4.15e-19
C5340 DVDD.n630 DGND 0.00105f
C5341 DVDD.t353 DGND 2.06e-19
C5342 DVDD.t355 DGND 1.62e-19
C5343 DVDD.n631 DGND 3.98e-19
C5344 DVDD.n632 DGND 8.64e-19
C5345 DVDD.n633 DGND 0.001598f
C5346 DVDD.n634 DGND 2.3e-19
C5347 DVDD.n635 DGND 0.001171f
C5348 DVDD.n636 DGND 0.00105f
C5349 DVDD.t397 DGND 0.001428f
C5350 DVDD.n637 DGND 0.001662f
C5351 DVDD.n638 DGND 0.001415f
C5352 DVDD.t181 DGND 5.49e-19
C5353 DVDD.n639 DGND 0.001052f
C5354 DVDD.n640 DGND 4.15e-19
C5355 DVDD.n641 DGND 0.001377f
C5356 DVDD.n642 DGND 0.00105f
C5357 DVDD.t86 DGND 3.58e-19
C5358 DVDD.t105 DGND 3.58e-19
C5359 DVDD.n643 DGND 7.77e-19
C5360 DVDD.n644 DGND 3.75e-19
C5361 DVDD.n645 DGND 0.00105f
C5362 DVDD.t207 DGND 7.66e-19
C5363 DVDD.n646 DGND 0.001178f
C5364 DVDD.n647 DGND 0.001641f
C5365 DVDD.t205 DGND 0.001258f
C5366 DVDD.n648 DGND 7.9e-19
C5367 DVDD.n649 DGND 0.003071f
C5368 DVDD.n650 DGND 3.39e-19
C5369 DVDD.n651 DGND 0.00105f
C5370 DVDD.n652 DGND 0.00105f
C5371 DVDD.n653 DGND 2.62e-19
C5372 DVDD.n654 DGND 4.15e-19
C5373 DVDD.n655 DGND 0.00105f
C5374 DVDD.n656 DGND 0.00105f
C5375 DVDD.n657 DGND 2.12e-19
C5376 DVDD.n658 DGND 9.14e-19
C5377 DVDD.n659 DGND 4.99e-19
C5378 DVDD.n660 DGND 0.00105f
C5379 DVDD.n661 DGND 0.00105f
C5380 DVDD.n662 DGND 2.23e-19
C5381 DVDD.t295 DGND 1.51e-19
C5382 DVDD.t114 DGND 1.51e-19
C5383 DVDD.n663 DGND 3.12e-19
C5384 DVDD.n664 DGND 9.76e-19
C5385 DVDD.n665 DGND 2.5e-19
C5386 DVDD.n666 DGND 2.32e-19
C5387 DVDD.n667 DGND 0.001552f
C5388 DVDD.n668 DGND 0.001377f
C5389 DVDD.n669 DGND 3.59e-19
C5390 DVDD.n670 DGND 0.00105f
C5391 DVDD.n671 DGND 0.00105f
C5392 DVDD.t334 DGND 1.51e-19
C5393 DVDD.t133 DGND 1.51e-19
C5394 DVDD.n672 DGND 3.12e-19
C5395 DVDD.n673 DGND 0.001184f
C5396 DVDD.n674 DGND 2.78e-19
C5397 DVDD.n675 DGND 4.15e-19
C5398 DVDD.n676 DGND 0.00137f
C5399 DVDD.n677 DGND 0.001377f
C5400 DVDD.n678 DGND 3.99e-19
C5401 DVDD.n679 DGND 0.00105f
C5402 DVDD.n680 DGND 0.00105f
C5403 DVDD.n681 DGND 3.86e-19
C5404 DVDD.t55 DGND 7.6e-19
C5405 DVDD.n682 DGND 0.001385f
C5406 DVDD.n683 DGND 0.00105f
C5407 DVDD.n684 DGND 0.00105f
C5408 DVDD.n685 DGND 4.15e-19
C5409 DVDD.n686 DGND 4.15e-19
C5410 DVDD.n687 DGND 4.15e-19
C5411 DVDD.n688 DGND 0.001598f
C5412 DVDD.n689 DGND 0.001253f
C5413 DVDD.n690 DGND 0.001919f
C5414 DVDD.n691 DGND 0.005545f
C5415 DVDD.t390 DGND 0.01244f
C5416 DVDD.t43 DGND 0.01129f
C5417 DVDD.t54 DGND 0.003067f
C5418 DVDD.t352 DGND 0.00409f
C5419 DVDD.t296 DGND 0.00409f
C5420 DVDD.t354 DGND 0.003067f
C5421 DVDD.t130 DGND 0.006263f
C5422 DVDD.t214 DGND 0.007882f
C5423 DVDD.t333 DGND 0.00737f
C5424 DVDD.t132 DGND 0.004899f
C5425 DVDD.t396 DGND 0.003579f
C5426 DVDD.t180 DGND 0.010267f
C5427 DVDD.t294 DGND 0.011332f
C5428 DVDD.t476 DGND 0.003579f
C5429 DVDD.t113 DGND 0.003579f
C5430 DVDD.t85 DGND 0.003579f
C5431 DVDD.t131 DGND 0.003579f
C5432 DVDD.t104 DGND 0.003579f
C5433 DVDD.t19 DGND 0.003579f
C5434 DVDD.t204 DGND 0.003834f
C5435 DVDD.t206 DGND 0.008009f
C5436 DVDD.t434 DGND 0.017254f
C5437 DVDD.t436 DGND 0.011503f
C5438 DVDD.t42 DGND 0.014144f
C5439 DVDD.t520 DGND 0.00605f
C5440 DVDD.t423 DGND 0.005794f
C5441 DVDD.t408 DGND 0.003579f
C5442 DVDD.t217 DGND 0.003579f
C5443 DVDD.t108 DGND 0.003579f
C5444 DVDD.t465 DGND 0.003579f
C5445 DVDD.t184 DGND 0.003579f
C5446 DVDD.t182 DGND 0.003579f
C5447 DVDD.t381 DGND 0.008009f
C5448 DVDD.t157 DGND 0.009628f
C5449 DVDD.t218 DGND 0.007157f
C5450 DVDD.t499 DGND 0.003962f
C5451 DVDD.t373 DGND 0.003792f
C5452 DVDD.t316 DGND 0.007498f
C5453 DVDD.t221 DGND 0.007157f
C5454 DVDD.t406 DGND 0.005411f
C5455 DVDD.n692 DGND 0.005247f
C5456 DVDD.n693 DGND 0.001919f
C5457 DVDD.n694 DGND 0.001892f
C5458 DVDD.n695 DGND 0.00105f
C5459 DVDD.n696 DGND 3.86e-19
C5460 DVDD.n697 DGND 4.15e-19
C5461 DVDD.n698 DGND 0.001735f
C5462 DVDD.n699 DGND 0.001233f
C5463 DVDD.n700 DGND 0.001171f
C5464 DVDD.t374 DGND 0.001428f
C5465 DVDD.n701 DGND 0.001662f
C5466 DVDD.n702 DGND 3.59e-19
C5467 DVDD.n703 DGND 0.00105f
C5468 DVDD.n704 DGND 0.00105f
C5469 DVDD.n705 DGND 2.78e-19
C5470 DVDD.n706 DGND 0.001184f
C5471 DVDD.n707 DGND 2.3e-19
C5472 DVDD.n708 DGND 0.001918f
C5473 DVDD.n709 DGND 4.07e-19
C5474 DVDD.n710 DGND 0.002427f
C5475 DVDD.n711 DGND 2.32e-19
C5476 DVDD.n712 DGND 2.5e-19
C5477 DVDD.n713 DGND 9.76e-19
C5478 DVDD.n714 DGND 4.15e-19
C5479 DVDD.n715 DGND 2.23e-19
C5480 DVDD.n716 DGND 0.0021f
C5481 DVDD.n717 DGND 2.12e-19
C5482 DVDD.n718 DGND 3.75e-19
C5483 DVDD.n719 DGND 7.9e-19
C5484 DVDD.n720 DGND 3.39e-19
C5485 DVDD.n721 DGND 0.0021f
C5486 DVDD.n722 DGND 0.0021f
C5487 DVDD.n723 DGND 2.62e-19
C5488 DVDD.n724 DGND 0.001178f
C5489 DVDD.n725 DGND 0.002811f
C5490 DVDD.n726 DGND 0.012547f
C5491 DVDD.n727 DGND 0.018412f
C5492 DVDD.n728 DGND 0.002811f
C5493 DVDD.t318 DGND 7.66e-19
C5494 DVDD.n729 DGND 0.001178f
C5495 DVDD.n730 DGND 2.62e-19
C5496 DVDD.n731 DGND 0.0021f
C5497 DVDD.n732 DGND 0.0021f
C5498 DVDD.n733 DGND 3.39e-19
C5499 DVDD.n734 DGND 7.9e-19
C5500 DVDD.n735 DGND 3.75e-19
C5501 DVDD.n736 DGND 2.12e-19
C5502 DVDD.n737 DGND 0.0021f
C5503 DVDD.n738 DGND 0.0021f
C5504 DVDD.n739 DGND 2.5e-19
C5505 DVDD.n740 DGND 2.32e-19
C5506 DVDD.t364 DGND 5.49e-19
C5507 DVDD.n741 DGND 0.001052f
C5508 DVDD.n742 DGND 2.3e-19
C5509 DVDD.n743 DGND 0.001918f
C5510 DVDD.n744 DGND 0.001377f
C5511 DVDD.n745 DGND 3.59e-19
C5512 DVDD.n746 DGND 0.00105f
C5513 DVDD.n747 DGND 0.00105f
C5514 DVDD.n748 DGND 2.78e-19
C5515 DVDD.n749 DGND 4.15e-19
C5516 DVDD.n750 DGND 0.001233f
C5517 DVDD.n751 DGND 0.001735f
C5518 DVDD.t304 DGND 0.004644f
C5519 DVDD.t336 DGND 0.003579f
C5520 DVDD.t134 DGND 0.00409f
C5521 DVDD.t187 DGND 0.00409f
C5522 DVDD.t319 DGND 0.003067f
C5523 DVDD.t251 DGND 0.004644f
C5524 DVDD.t398 DGND 0.007882f
C5525 DVDD.t151 DGND 0.00737f
C5526 DVDD.t252 DGND 0.004899f
C5527 DVDD.t238 DGND 0.003579f
C5528 DVDD.t382 DGND 0.010267f
C5529 DVDD.t324 DGND 0.011332f
C5530 DVDD.t225 DGND 0.003579f
C5531 DVDD.t176 DGND 0.003579f
C5532 DVDD.t417 DGND 0.003579f
C5533 DVDD.t254 DGND 0.003579f
C5534 DVDD.t424 DGND 0.003579f
C5535 DVDD.t165 DGND 0.003579f
C5536 DVDD.t361 DGND 0.003834f
C5537 DVDD.t73 DGND 0.008009f
C5538 DVDD.t186 DGND 0.017254f
C5539 DVDD.t38 DGND 0.011503f
C5540 DVDD.t531 DGND 0.014144f
C5541 DVDD.t317 DGND 0.00605f
C5542 DVDD.t435 DGND 0.005794f
C5543 DVDD.t367 DGND 0.003579f
C5544 DVDD.t0 DGND 0.003579f
C5545 DVDD.t287 DGND 0.003579f
C5546 DVDD.t458 DGND 0.003579f
C5547 DVDD.t96 DGND 0.003579f
C5548 DVDD.t117 DGND 0.003579f
C5549 DVDD.t6 DGND 0.008009f
C5550 DVDD.t363 DGND 0.009628f
C5551 DVDD.t1 DGND 0.007157f
C5552 DVDD.t106 DGND 0.003962f
C5553 DVDD.t78 DGND 0.003792f
C5554 DVDD.t375 DGND 0.007498f
C5555 DVDD.t3 DGND 0.007157f
C5556 DVDD.t12 DGND 0.005411f
C5557 DVDD.n752 DGND 0.005247f
C5558 DVDD.n753 DGND 0.001919f
C5559 DVDD.n754 DGND 0.001253f
C5560 DVDD.n755 DGND 0.00105f
C5561 DVDD.n756 DGND 3.86e-19
C5562 DVDD.t39 DGND 7.6e-19
C5563 DVDD.n757 DGND 0.001385f
C5564 DVDD.n758 DGND 0.002659f
C5565 DVDD.n759 DGND 0.003071f
C5566 DVDD.n760 DGND 3.39e-19
C5567 DVDD.n761 DGND 0.00105f
C5568 DVDD.n762 DGND 0.00105f
C5569 DVDD.n763 DGND 2.62e-19
C5570 DVDD.n764 DGND 4.15e-19
C5571 DVDD.n765 DGND 0.00105f
C5572 DVDD.n766 DGND 0.00105f
C5573 DVDD.n767 DGND 2.12e-19
C5574 DVDD.n768 DGND 9.14e-19
C5575 DVDD.n769 DGND 4.99e-19
C5576 DVDD.n770 DGND 0.00105f
C5577 DVDD.n771 DGND 0.00105f
C5578 DVDD.n772 DGND 2.23e-19
C5579 DVDD.t325 DGND 1.51e-19
C5580 DVDD.t177 DGND 1.51e-19
C5581 DVDD.n773 DGND 3.12e-19
C5582 DVDD.n774 DGND 9.76e-19
C5583 DVDD.n775 DGND 2.5e-19
C5584 DVDD.n776 DGND 2.32e-19
C5585 DVDD.n777 DGND 0.001552f
C5586 DVDD.n778 DGND 0.001377f
C5587 DVDD.n779 DGND 3.59e-19
C5588 DVDD.n780 DGND 0.00105f
C5589 DVDD.n781 DGND 0.00105f
C5590 DVDD.t152 DGND 1.51e-19
C5591 DVDD.t253 DGND 1.51e-19
C5592 DVDD.n782 DGND 3.12e-19
C5593 DVDD.n783 DGND 0.001184f
C5594 DVDD.n784 DGND 2.78e-19
C5595 DVDD.n785 DGND 4.15e-19
C5596 DVDD.n786 DGND 0.00137f
C5597 DVDD.n787 DGND 0.00105f
C5598 DVDD.n788 DGND 0.001517f
C5599 DVDD.n789 DGND 3.45e-19
C5600 DVDD.n790 DGND 0.00105f
C5601 DVDD.n791 DGND 0.00105f
C5602 DVDD.n792 DGND 3.86e-19
C5603 DVDD.t337 DGND 7.6e-19
C5604 DVDD.n793 DGND 0.001385f
C5605 DVDD.n794 DGND 0.00105f
C5606 DVDD.n795 DGND 0.00105f
C5607 DVDD.n796 DGND 3.41e-19
C5608 DVDD.n797 DGND 0.001838f
C5609 DVDD.n798 DGND 0.001918f
C5610 DVDD.n799 DGND 0.00212f
C5611 DVDD.n800 DGND 0.001919f
C5612 DVDD.n801 DGND 0.014407f
C5613 DVDD.t302 DGND 0.020888f
C5614 DVDD.n802 DGND 0.015646f
C5615 DVDD.t128 DGND 0.013936f
C5616 DVDD.t249 DGND 0.004644f
C5617 DVDD.t40 DGND 0.003579f
C5618 DVDD.t399 DGND 0.00409f
C5619 DVDD.t393 DGND 0.00409f
C5620 DVDD.t450 DGND 0.003067f
C5621 DVDD.t127 DGND 0.004644f
C5622 DVDD.t110 DGND 0.007882f
C5623 DVDD.t255 DGND 0.00737f
C5624 DVDD.t124 DGND 0.004899f
C5625 DVDD.t350 DGND 0.003579f
C5626 DVDD.t163 DGND 0.010267f
C5627 DVDD.t178 DGND 0.011332f
C5628 DVDD.t501 DGND 0.003579f
C5629 DVDD.t474 DGND 0.003579f
C5630 DVDD.t153 DGND 0.003579f
C5631 DVDD.t126 DGND 0.003579f
C5632 DVDD.t83 DGND 0.003579f
C5633 DVDD.t247 DGND 0.003579f
C5634 DVDD.t517 DGND 0.003834f
C5635 DVDD.t228 DGND 0.008009f
C5636 DVDD.t137 DGND 0.017254f
C5637 DVDD.t344 DGND 0.011503f
C5638 DVDD.n803 DGND 0.005247f
C5639 DVDD.n804 DGND 0.001919f
C5640 DVDD.n805 DGND 0.001253f
C5641 DVDD.n806 DGND 0.001735f
C5642 DVDD.n807 DGND 0.001233f
C5643 DVDD.n808 DGND 4.15e-19
C5644 DVDD.n809 DGND 2.78e-19
C5645 DVDD.n810 DGND 0.00105f
C5646 DVDD.n811 DGND 0.00105f
C5647 DVDD.n812 DGND 3.59e-19
C5648 DVDD.n813 DGND 0.001377f
C5649 DVDD.n814 DGND 0.001918f
C5650 DVDD.n815 DGND 2.3e-19
C5651 DVDD.t534 DGND 5.49e-19
C5652 DVDD.n816 DGND 0.001052f
C5653 DVDD.n817 DGND 2.32e-19
C5654 DVDD.n818 DGND 2.5e-19
C5655 DVDD.n819 DGND 0.0021f
C5656 DVDD.n820 DGND 4.07e-19
C5657 DVDD.n821 DGND 0.001006f
C5658 DVDD.n822 DGND 2.12e-19
C5659 DVDD.n823 DGND 3.75e-19
C5660 DVDD.n824 DGND 0.0021f
C5661 DVDD.n825 DGND 0.0021f
C5662 DVDD.n826 DGND 0.0021f
C5663 DVDD.n827 DGND 4.12e-19
C5664 DVDD.n828 DGND 0.002811f
C5665 DVDD.n829 DGND 0.018412f
C5666 DVDD.n830 DGND 0.002178f
C5667 DVDD.n831 DGND 0.001178f
C5668 DVDD.n832 DGND 2.62e-19
C5669 DVDD.n833 DGND 4.15e-19
C5670 DVDD.n834 DGND 0.001172f
C5671 DVDD.n835 DGND 0.001172f
C5672 DVDD.n836 DGND 0.001172f
C5673 DVDD.n837 DGND 2.23e-19
C5674 DVDD.n838 DGND 9.76e-19
C5675 DVDD.n839 DGND 2.5e-19
C5676 DVDD.n840 DGND 2.32e-19
C5677 DVDD.n841 DGND 0.001172f
C5678 DVDD.n842 DGND 0.001172f
C5679 DVDD.n843 DGND 2.3e-19
C5680 DVDD.n844 DGND 0.001184f
C5681 DVDD.n845 DGND 2.78e-19
C5682 DVDD.n846 DGND 0.001172f
C5683 DVDD.n847 DGND 0.001172f
C5684 DVDD.n848 DGND 0.001172f
C5685 DVDD.n849 DGND 4.15e-19
C5686 DVDD.n850 DGND 3.86e-19
C5687 DVDD.n851 DGND 0.001385f
C5688 DVDD.n852 DGND 0.002231f
C5689 DVDD.n853 DGND 0.002282f
C5690 DVDD.n854 DGND 0.001178f
C5691 DVDD.n855 DGND 2.62e-19
C5692 DVDD.n856 DGND 4.15e-19
C5693 DVDD.n857 DGND 0.001172f
C5694 DVDD.n858 DGND 0.001172f
C5695 DVDD.n859 DGND 0.001172f
C5696 DVDD.n860 DGND 2.23e-19
C5697 DVDD.n861 DGND 9.76e-19
C5698 DVDD.n862 DGND 2.5e-19
C5699 DVDD.n863 DGND 2.32e-19
C5700 DVDD.n864 DGND 0.001172f
C5701 DVDD.n865 DGND 0.001172f
C5702 DVDD.n866 DGND 2.3e-19
C5703 DVDD.n867 DGND 0.001184f
C5704 DVDD.n868 DGND 2.78e-19
C5705 DVDD.n869 DGND 0.001172f
C5706 DVDD.n870 DGND 0.001172f
C5707 DVDD.n871 DGND 0.001172f
C5708 DVDD.n872 DGND 4.15e-19
C5709 DVDD.n873 DGND 3.86e-19
C5710 DVDD.n874 DGND 0.001385f
C5711 DVDD.n875 DGND 0.002623f
C5712 DVDD.t308 DGND 0.010097f
C5713 DVDD.t248 DGND 0.003706f
C5714 DVDD.t410 DGND 0.003579f
C5715 DVDD.t160 DGND 0.003579f
C5716 DVDD.t16 DGND 0.005794f
C5717 DVDD.t155 DGND 0.005794f
C5718 DVDD.t379 DGND 0.003579f
C5719 DVDD.t310 DGND 0.003685f
C5720 DVDD.t346 DGND 0.003941f
C5721 DVDD.t150 DGND 0.003579f
C5722 DVDD.t123 DGND 0.003579f
C5723 DVDD.t8 DGND 0.010672f
C5724 DVDD.t174 DGND 0.010544f
C5725 DVDD.t75 DGND 0.003706f
C5726 DVDD.t268 DGND 0.003579f
C5727 DVDD.t35 DGND 0.003579f
C5728 DVDD.t244 DGND 0.005794f
C5729 DVDD.t208 DGND 0.005794f
C5730 DVDD.t266 DGND 0.003579f
C5731 DVDD.t504 DGND 0.003685f
C5732 DVDD.t349 DGND 0.003941f
C5733 DVDD.t265 DGND 0.003579f
C5734 DVDD.t467 DGND 0.003579f
C5735 DVDD.t33 DGND 0.01205f
C5736 DVDD.n876 DGND 0.018801f
C5737 DVDD.t94 DGND 0.010097f
C5738 DVDD.t404 DGND 0.003706f
C5739 DVDD.t496 DGND 0.003579f
C5740 DVDD.t536 DGND 0.003579f
C5741 DVDD.t68 DGND 0.005794f
C5742 DVDD.t70 DGND 0.005794f
C5743 DVDD.t497 DGND 0.003579f
C5744 DVDD.t430 DGND 0.003685f
C5745 DVDD.t80 DGND 0.003941f
C5746 DVDD.t480 DGND 0.003579f
C5747 DVDD.t405 DGND 0.003579f
C5748 DVDD.t432 DGND 0.010672f
C5749 DVDD.t428 DGND 0.010544f
C5750 DVDD.t535 DGND 0.003706f
C5751 DVDD.t145 DGND 0.003579f
C5752 DVDD.t421 DGND 0.003579f
C5753 DVDD.t369 DGND 0.005794f
C5754 DVDD.t477 DGND 0.005794f
C5755 DVDD.t142 DGND 0.003579f
C5756 DVDD.t426 DGND 0.003685f
C5757 DVDD.t240 DGND 0.003941f
C5758 DVDD.t144 DGND 0.003579f
C5759 DVDD.t291 DGND 0.003579f
C5760 DVDD.t419 DGND 0.01205f
C5761 DVDD.n877 DGND 0.018801f
C5762 DVDD.n878 DGND 0.002623f
C5763 DVDD.t420 DGND 7.6e-19
C5764 DVDD.n879 DGND 0.001385f
C5765 DVDD.n880 DGND 3.86e-19
C5766 DVDD.n881 DGND 4.15e-19
C5767 DVDD.n882 DGND 0.001172f
C5768 DVDD.n883 DGND 0.001172f
C5769 DVDD.n884 DGND 0.001172f
C5770 DVDD.n885 DGND 2.78e-19
C5771 DVDD.n886 DGND 0.001184f
C5772 DVDD.n887 DGND 2.3e-19
C5773 DVDD.n888 DGND 0.001172f
C5774 DVDD.n889 DGND 0.001172f
C5775 DVDD.n890 DGND 2.32e-19
C5776 DVDD.n891 DGND 2.5e-19
C5777 DVDD.n892 DGND 9.76e-19
C5778 DVDD.n893 DGND 2.23e-19
C5779 DVDD.n894 DGND 0.001172f
C5780 DVDD.n895 DGND 0.001172f
C5781 DVDD.n896 DGND 0.001172f
C5782 DVDD.n897 DGND 4.15e-19
C5783 DVDD.n898 DGND 2.62e-19
C5784 DVDD.n899 DGND 0.001178f
C5785 DVDD.n900 DGND 0.002282f
C5786 DVDD.t433 DGND 7.6e-19
C5787 DVDD.n901 DGND 0.001385f
C5788 DVDD.n902 DGND 0.002231f
C5789 DVDD.n903 DGND 0.00143f
C5790 DVDD.n904 DGND 0.001172f
C5791 DVDD.n905 DGND 4.15e-19
C5792 DVDD.n906 DGND 4.15e-19
C5793 DVDD.n907 DGND 2.78e-19
C5794 DVDD.n908 DGND 0.001172f
C5795 DVDD.n909 DGND 0.001172f
C5796 DVDD.n910 DGND 0.001172f
C5797 DVDD.n911 DGND 2.3e-19
C5798 DVDD.n912 DGND 0.001052f
C5799 DVDD.n913 DGND 2.32e-19
C5800 DVDD.t69 DGND 1.51e-19
C5801 DVDD.t537 DGND 1.51e-19
C5802 DVDD.n914 DGND 3.12e-19
C5803 DVDD.n915 DGND 9.76e-19
C5804 DVDD.n916 DGND 2.5e-19
C5805 DVDD.n917 DGND 0.001172f
C5806 DVDD.n918 DGND 0.001172f
C5807 DVDD.n919 DGND 0.001172f
C5808 DVDD.n920 DGND 4.15e-19
C5809 DVDD.n921 DGND 4.15e-19
C5810 DVDD.t95 DGND 7.66e-19
C5811 DVDD.n922 DGND 0.001178f
C5812 DVDD.n923 DGND 2.62e-19
C5813 DVDD.n924 DGND 7.13e-19
.ends

