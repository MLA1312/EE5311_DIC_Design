** sch_path: /home/EE23B038/ee5311/tutorial_3/tutorial_3_1c.sch
**.subckt tutorial_3_1c
XM2 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vin1 Vin GND 1.8
Vdd1 VDD GND 1.8
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.control
let vds = 0.2
set vtccache = ( )
set idscache = ( )
let index = 1
let N = 10
let imax = vector(N)
let vdscache = vector(N)
while index le N
    alter Vdd1 $&vds
    dc Vin1 0 $&vds 0.01
    set vtccache = ( $vtccache dc{$&index}.v(Vout) )
    set idscache = ( $idscache dc{$&index}.i(Vdd1) )
    let imax[index - 1] = abs(vecmin(dc{$&index}.i(Vdd1)))
    let vdscache[index - 1] = vds
    let vds = vds + 0.2
    let index = index + 1
end
plot $vtccache
plot $idscache
plot imax vs vdscache
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
