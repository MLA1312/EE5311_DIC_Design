** sch_path: /home/EE23B038/ee5311/tutorial_4/tutorial_4_2a.sch
**.subckt tutorial_4_2a
x1 net1 Vout inv
x2 net2 net1 inv
x3 net3 net2 inv
x4 net4 net3 inv
x5 net5 net4 inv
x6 net6 net5 inv
x7 Vout net6 inv
Vdd1 VDD GND 1.8
**** begin user architecture code


.ic v(Vout) = 0
.param width_p = 0.84
.control
tran 0.001n 1n
plot v(Vout)
meas tran period trig v(Vout) val=0.9 rise=1 targ v(Vout) val=0.9 rise=2
let freq = 1/ $&period
echo freq: $&freq
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  /home/EE23B038/ee5311/tutorial_4/inv.sym # of pins=2
** sym_path: /home/EE23B038/ee5311/tutorial_4/inv.sym
** sch_path: /home/EE23B038/ee5311/tutorial_4/inv.sch
.subckt inv out in
*.ipin in
*.opin out
XM1 out in GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W={width_p} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
