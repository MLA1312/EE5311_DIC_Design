** sch_path: /home/EE23B038/ee5311/tutorial_2/tutorial_2_2b.sch
**.subckt tutorial_2_2b
XM2 net3 net2 net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdd1 net1 GND 1.8
Vin1 net2 GND 1.8
Vdr1 net3 GND 1.8
**** begin user architecture code


.control
let Vg = 1.2
let mu = 0.009
let WbyL = 0.42/0.15
let Cox = 0.00816
let Vth = 0.7
let vsat = 3e4
let lambdap = 0.2
let EcL = 2*vsat* 0.15e-6/mu
repeat 4
   alter Vin1 $&Vg
   dc Vdr1 1.8 0 -0.02
   let Vsd = 1.8 - "v-sweep"
   let Vsg = 1.8 - Vg
   let Vsd1 = min(Vsg - Vth, Vsd)
   let Vgt = max(Vsg - Vth, 0)
   let Vsd_min = min(Vsd1, EcL*Vgt/(EcL+Vgt))
   let idfit = mu*Cox*WbyL*EcL*(Vsg - Vth - Vsd_min/2)*Vsd_min*(1 + lambdap * Vsd)/(Vsd_min + EcL)
   let Vg = Vg - 0.4
end
plot dc1.I(Vdr1) dc2.I(Vdr1) dc3.I(Vdr1) dc4.I(Vdr1) dc1.idfit dc2.idfit dc3.idfit dc4.idfit
set filetype=ascii
wrdata pmos_ids_vds.txt dc1.I(Vdr1) dc2.I(Vdr1) dc3.I(Vdr1) dc4.I(Vdr1) dc1.idfit dc2.idfit dc3.idfit dc4.idfit
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
