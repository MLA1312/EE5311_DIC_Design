* NGSPICE file created from ring_osc.ext - technology: sky130A
.subckt ring_osc DVDD val DGND
X0 a_973_41# a_493_41# DGND.t11 DGND.t10 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 a_1453_41# a_973_41# DVDD.t13 DVDD.t12 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X2 a_1933_41# a_1453_41# DVDD.t1 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X3 a_1453_41# a_973_41# DGND.t13 DGND.t12 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X4 a_2413_41# a_1933_41# DGND.t7 DGND.t6 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X5 a_13_41# val.t2 DGND.t9 DGND.t8 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X6 a_2413_41# a_1933_41# DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X7 val.t1 a_2413_41# DVDD.t3 DVDD.t2 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X8 a_493_41# a_13_41# DGND.t5 DGND.t4 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X9 a_1933_41# a_1453_41# DGND.t1 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X10 val.t0 a_2413_41# DGND.t3 DGND.t2 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X11 a_13_41# val.t3 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X12 a_493_41# a_13_41# DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X13 a_973_41# a_493_41# DVDD.t11 DVDD.t10 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
R0 DGND.t2 DGND.n2 4634.22
R1 DGND.n3 DGND.t2 3417.48
R2 DGND.t6 DGND.n3 3417.48
R3 DGND.n15 DGND.t6 3417.48
R4 DGND.n15 DGND.t0 3417.48
R5 DGND.t0 DGND.n14 3417.48
R6 DGND.n14 DGND.t12 3417.48
R7 DGND.n10 DGND.t12 3417.48
R8 DGND.n10 DGND.t10 3417.48
R9 DGND.t10 DGND.n9 3417.48
R10 DGND.n9 DGND.t4 3417.48
R11 DGND.n5 DGND.t4 3417.48
R12 DGND.n5 DGND.t8 3417.48
R13 DGND.n6 DGND.n5 1216.38
R14 DGND.n9 DGND.n8 1216.38
R15 DGND.n11 DGND.n10 1216.38
R16 DGND.n14 DGND.n13 1216.38
R17 DGND.n16 DGND.n15 1216.38
R18 DGND.n3 DGND.n0 1216.38
R19 DGND.n6 DGND.t9 276.111
R20 DGND.n7 DGND.t5 275.74
R21 DGND.n4 DGND.t11 275.74
R22 DGND.n12 DGND.t13 275.74
R23 DGND.n1 DGND.t1 275.74
R24 DGND.n17 DGND.t7 275.74
R25 DGND.n2 DGND.t3 275.74
R26 DGND.n16 DGND.n1 0.371594
R27 DGND.n13 DGND.n12 0.371594
R28 DGND.n11 DGND.n4 0.371594
R29 DGND.n8 DGND.n7 0.371594
R30 DGND.n2 DGND.n0 0.254406
R31 DGND.n17 DGND.n16 0.254406
R32 DGND.n13 DGND.n1 0.254406
R33 DGND.n12 DGND.n11 0.254406
R34 DGND.n8 DGND.n4 0.254406
R35 DGND.n7 DGND.n6 0.254406
R36 DGND DGND.n0 0.237479
R37 DGND DGND.n17 0.134615
R38 DVDD.t2 DVDD.n2 942.977
R39 DVDD.n3 DVDD.t2 703.705
R40 DVDD.n3 DVDD.t8 703.705
R41 DVDD.n7 DVDD.t8 703.705
R42 DVDD.t0 DVDD.n7 703.705
R43 DVDD.n16 DVDD.t0 703.705
R44 DVDD.n16 DVDD.t12 703.705
R45 DVDD.t12 DVDD.n15 703.705
R46 DVDD.n15 DVDD.t10 703.705
R47 DVDD.n11 DVDD.t10 703.705
R48 DVDD.n11 DVDD.t4 703.705
R49 DVDD.t4 DVDD.n10 703.705
R50 DVDD.n10 DVDD.t6 703.705
R51 DVDD.n9 DVDD.t7 398.221
R52 DVDD.n8 DVDD.t5 397.849
R53 DVDD.n13 DVDD.t11 397.849
R54 DVDD.n1 DVDD.t13 397.849
R55 DVDD.n0 DVDD.t1 397.849
R56 DVDD.n5 DVDD.t9 397.849
R57 DVDD.n2 DVDD.t3 397.849
R58 DVDD.n4 DVDD.n3 238.904
R59 DVDD.n7 DVDD.n6 238.904
R60 DVDD.n17 DVDD.n16 238.904
R61 DVDD.n15 DVDD.n14 238.904
R62 DVDD.n12 DVDD.n11 238.904
R63 DVDD.n10 DVDD.n9 238.904
R64 DVDD.n5 DVDD.n4 0.371594
R65 DVDD.n6 DVDD.n0 0.371594
R66 DVDD.n17 DVDD.n1 0.371594
R67 DVDD.n14 DVDD.n13 0.371594
R68 DVDD.n12 DVDD.n8 0.371594
R69 DVDD.n4 DVDD.n2 0.254406
R70 DVDD.n6 DVDD.n5 0.254406
R71 DVDD.n14 DVDD.n1 0.254406
R72 DVDD.n13 DVDD.n12 0.254406
R73 DVDD.n9 DVDD.n8 0.254406
R74 DVDD DVDD.n17 0.146333
R75 DVDD DVDD.n0 0.108573
R76 val.n0 val.t1 407.534
R77 val.n0 val.t0 271.118
R78 val.n1 val.t3 260.779
R79 val.n1 val.t2 177.232
R80 val val.n1 168.183
R81 val val.n0 9.3167
C0 a_493_41# a_13_41# 0.059446f
C1 a_973_41# val 0.09771f
C2 DVDD a_13_41# 0.272156f
C3 a_1453_41# DVDD 0.278798f
C4 a_493_41# val 0.09771f
C5 DVDD a_1933_41# 0.278798f
C6 DVDD val 0.902631f
C7 val a_13_41# 0.150352f
C8 a_1453_41# a_1933_41# 0.059446f
C9 a_1453_41# val 0.09771f
C10 a_2413_41# DVDD 0.277024f
C11 val a_1933_41# 0.09771f
C12 a_973_41# a_493_41# 0.059446f
C13 a_2413_41# a_1933_41# 0.059446f
C14 a_973_41# DVDD 0.278798f
C15 a_2413_41# val 0.144679f
C16 a_973_41# a_1453_41# 0.059446f
C17 a_493_41# DVDD 0.278798f
C18 val DGND 1.12115f
C19 DVDD DGND 4.21912f
C20 a_2413_41# DGND 0.395776f
C21 a_1933_41# DGND 0.384637f
C22 a_1453_41# DGND 0.384637f
C23 a_973_41# DGND 0.384637f
C24 a_493_41# DGND 0.384637f
C25 a_13_41# DGND 0.400555f
.ends
