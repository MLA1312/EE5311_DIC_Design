* NGSPICE file created from fa16.ext - technology: sky130A

.subckt fa16 DGND DVDD B4 A4 A5 B5 B6 A6 A7 B7 A8 B8 A9 B9 S15 B10 A10 A11 B11 B12
+ A12 A13 B13 B14 A14 A15 B15 B0 A0 A1 B1 B2 A2 A3 B3 Cin
X0 a_4691_n3974# A11 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_5402_n3546# a_4204_n3054# a_5819_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_4691_n1494# A15 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_541_n828# A2 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 DVDD a_1201_n3054# a_2273_n2734# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X5 a_5288_n828# B14 a_5192_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 DGND B9 a_4363_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_4697_n2434# B9 a_3946_n2306# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_894_n1194# a_143_n1036# a_798_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 DGND A10 a_5456_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X10 a_894_n3674# a_143_n3516# a_798_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 DGND A14 a_5456_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X12 DVDD A2 a_n41_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_n131_n574# a_n71_n600# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X14 a_1467_46# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X15 a_4691_n1814# A15 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 DVDD A6 a_185_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_11_n1194# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X18 a_3874_n3700# a_5402_n3546# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_11_n3674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X20 a_3874_n1220# a_5402_n1066# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_5819_n2068# A8 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 DVDD a_3861_n3080# a_3322_n4062# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X23 a_147_n1494# B2 a_n131_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X24 a_147_n3974# B6 a_n131_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X25 a_315_n3054# A4 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 DGND B2 a_n71_n1840# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 DGND B6 a_n71_n4320# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_3832_46# B13 a_3736_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_3655_n1516# a_3322_n1582# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_966_n3674# B6 a_894_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 a_4523_n3054# B9 a_4441_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_2350_46# a_636_n574# a_2254_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_3874_20# a_5402_174# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X34 a_966_n1194# B2 a_894_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X35 DGND A11 a_4441_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 DGND A15 a_4441_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 a_3765_n3080# a_4441_n3054# a_4691_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X38 DVDD B10 a_5456_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 a_3736_n3308# A11 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X40 a_3874_n1220# a_5402_n1066# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X41 DVDD A13 a_4523_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X42 a_5192_n1194# A14 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X43 a_5192_n3674# A10 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X44 DVDD a_1557_n2434# a_143_n3516# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X45 a_2273_n254# a_1201_n1814# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 a_n71_n600# B0 a_315_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X47 DGND A7 a_1641_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X48 a_6153_n2068# B8 a_5402_n2306# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X49 a_n41_n1814# B2 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X50 DGND A3 a_1641_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X51 a_n41_n1814# a_n71_n1840# a_n131_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X52 a_1641_412# a_636_n574# a_1557_46# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X53 a_5819_n828# A14 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X54 a_n71_n1840# B2 a_315_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X55 a_3765_n3080# B9 a_4691_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X56 DVDD A15 a_4523_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X57 a_4697_n828# B15 a_3946_n1066# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X58 a_11_46# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X59 a_5360_n2434# a_2995_n4294# a_5288_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X60 a_541_n828# B2 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X61 DVDD A10 a_5855_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X62 DVDD A0 a_185_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X63 DVDD A13 a_4697_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X64 a_1641_n2434# a_636_n3054# a_1557_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 a_4000_n2068# a_3946_n2306# a_3904_n2434# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 DVDD B12 a_6023_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X67 a_894_n828# a_143_n1036# a_798_n1194# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_2422_n2434# B5 a_2350_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X69 a_185_n2068# B4 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X70 a_3655_n3996# a_3322_n4062# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 DVDD A10 a_6153_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X72 DVDD a_2908_n600# S15 DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X73 a_3655_n3996# a_3322_n4062# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X74 a_3655_n1516# a_3322_n1582# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X75 a_4000_46# a_3946_174# a_3904_46# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_1467_n1194# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X77 a_1467_n3674# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X78 a_5456_n3308# a_4204_n3054# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X79 DVDD A12 a_5456_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X80 a_1201_n3054# a_1261_n3080# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X81 DVDD a_636_n3054# a_1997_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X82 a_5402_n2306# a_2995_n4294# a_5819_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X83 a_101_n2434# B4 a_11_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X84 DGND B11 a_4363_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 DGND A0 a_185_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X86 a_4363_46# A13 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X87 DGND B15 a_4363_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X88 a_4697_n1194# B15 a_3946_n1066# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X89 a_4697_n3674# B11 a_3946_n3546# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 a_4697_412# B13 a_3946_174# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X91 DGND a_143_n2276# a_541_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X92 DVDD A15 a_4697_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X93 a_1557_n2434# B5 a_1467_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X94 DVDD a_3669_n342# a_3322_n1582# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 a_2790_n3928# a_1968_n4294# a_2569_n4255# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X96 a_798_n3674# a_101_n3674# a_541_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X97 a_1641_n2434# B5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X98 a_2790_n1448# a_1968_n1814# a_2569_n1775# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X99 DVDD A0 a_n41_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X100 a_4000_n2434# a_3874_n2460# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 DVDD A4 a_185_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X102 a_3543_n342# a_5773_n1814# a_6023_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X103 a_4697_46# B13 a_3946_174# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X104 a_6023_n254# A12 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 a_2908_n600# a_3874_n1220# a_3832_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X106 a_4363_n828# A15 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X107 a_3736_46# A13 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X108 a_185_412# Cin a_101_46# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X109 a_3832_n3308# B11 a_3736_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X110 a_1997_n3308# B7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X111 DGND A9 a_4697_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X112 a_315_n4294# A6 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X113 a_2254_46# a_1557_46# a_1997_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X114 DGND A5 a_1479_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X115 a_101_n1194# B2 a_11_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X116 DVDD A2 a_185_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X117 a_3946_n3546# a_3874_n3700# a_4363_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 a_4523_n4294# B11 a_4441_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X119 DGND a_5773_n574# a_3861_n600# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X120 a_3669_n2822# a_4441_n4294# a_4691_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X121 DVDD a_1557_n3674# a_1968_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X122 DVDD B8 a_5456_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 a_3736_n2068# A9 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X124 a_1557_46# B1 a_1467_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X125 DVDD A4 a_n41_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X126 DGND a_4441_n3054# a_3765_n3080# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X127 a_4204_n3054# a_3946_n2306# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X128 a_1997_n3308# A7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X129 a_4691_n3054# A9 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X130 a_3669_n2822# B11 a_4691_n3974# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X131 DGND a_5773_n3054# a_3861_n3080# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X132 a_3669_n342# B15 a_4691_n1494# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X133 a_2459_n254# a_1201_n574# a_2363_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X134 a_2254_n1194# a_1557_n1194# a_1997_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X135 DGND A9 a_4000_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X136 a_3946_174# a_3874_20# a_4363_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_5360_n1194# a_4204_n574# a_5288_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X138 a_5360_n3674# a_4204_n3054# a_5288_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X139 a_1641_n3674# a_636_n4294# a_1557_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 DVDD A6 a_966_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X141 DGND B1 a_1261_n600# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 a_3795_n254# a_3765_n600# a_3711_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X143 a_1641_n1194# a_636_n1814# a_1557_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X144 a_2422_n1194# B3 a_2350_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X145 a_2422_n3674# B7 a_2350_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X146 a_4000_46# a_3874_20# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X147 DVDD A8 a_6153_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X148 a_1479_n2734# B5 a_1201_n3054# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X149 a_4363_n3308# A11 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X150 a_3904_46# a_3874_20# a_3832_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X151 DVDD B15 a_4691_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X152 a_1467_412# A1 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X153 DGND A0 a_966_46# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X154 a_3874_n2460# a_5402_n2306# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X155 a_2422_46# B1 a_2350_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X156 a_5456_n2068# a_2995_n4294# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X157 a_1201_n1814# a_1261_n1840# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X158 a_1201_n4294# a_1261_n4320# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X159 a_966_n828# B2 a_894_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 a_n41_n3054# B4 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X161 a_n41_n3054# a_n71_n3080# a_n131_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X162 a_11_n828# A2 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X163 DVDD A14 a_5456_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X164 a_n71_n3080# B4 a_315_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X165 a_5855_n574# B12 a_5773_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X166 DVDD B15 a_4000_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 DVDD A10 a_5456_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X168 a_894_n3308# a_143_n3516# a_798_n3674# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X169 DVDD A9 a_4523_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 DVDD a_3861_n600# a_3322_n1582# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X171 DGND a_143_n3516# a_541_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X172 DGND a_143_n1036# a_541_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 a_6023_n2734# A8 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X174 a_6153_46# B12 a_5402_174# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X175 a_1557_n3674# B7 a_1467_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X176 a_1557_n1194# B3 a_1467_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X177 a_798_n2434# a_101_n2434# a_541_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X178 a_1641_n1194# B3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X179 a_1641_n3674# B7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 a_2497_n1775# a_2315_n1775# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X181 a_4000_n1194# a_3874_n1220# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X182 a_4000_n3674# a_3874_n3700# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X183 a_11_n3308# A6 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X184 a_541_412# B0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 a_541_n2434# B4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X186 a_1997_46# B1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X187 DVDD a_3226_n4062# a_3177_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X188 DGND A15 a_4697_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X189 DGND A11 a_4697_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X190 a_3832_n2068# B9 a_3736_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X191 a_1997_n2068# B5 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X192 DGND A1 a_1479_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X193 a_3627_n254# a_3543_n342# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X194 a_541_46# B0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X195 DGND A12 a_5456_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X196 a_147_n254# B0 a_n131_n574# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X197 DGND A3 a_1479_n1494# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X198 DGND A7 a_1479_n3974# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X199 a_966_n3308# B6 a_894_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X200 a_2254_n2434# a_1557_n2434# a_1997_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X201 a_2350_412# a_636_n574# a_2254_46# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X202 a_3946_n2306# a_3874_n2460# a_4363_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 a_5288_n2434# B8 a_5192_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X204 a_5192_n3308# A10 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X205 a_1641_n828# B3 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X206 a_2254_46# a_1557_46# a_1997_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X207 a_5360_46# a_3177_n4294# a_5288_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X208 a_894_46# Cin a_798_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X209 DVDD A6 a_n41_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X210 DGND a_4441_n4294# a_3669_n2822# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X211 DVDD A7 a_1641_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X212 a_2569_n1775# a_1968_n1814# a_2497_n1775# DVDD sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X213 a_3765_n600# a_4441_n574# a_4691_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X214 DGND a_4441_n1814# a_3669_n342# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X215 a_5192_46# A12 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X216 DGND A12 a_5773_n574# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X217 a_798_n1194# a_101_n1194# a_541_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X218 a_2497_n4255# a_2315_n4255# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_3434_n4026# a_3946_n3546# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X220 DGND B5 a_1261_n3080# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X221 a_1997_n2068# A5 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X222 a_3434_n1546# a_3946_n1066# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X223 a_4691_n4294# A11 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X224 DVDD A3 a_1291_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X225 a_3874_20# a_5402_174# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X226 DGND a_5773_n4294# a_3543_n2822# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X227 a_3861_n3080# a_5773_n3054# a_6023_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X228 DGND a_5773_n1814# a_3543_n342# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X229 a_4363_412# A13 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X230 DGND a_636_n574# a_1997_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X231 DGND A15 a_4000_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X232 DGND A11 a_4000_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X233 DVDD A4 a_966_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X234 DVDD A15 a_4000_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X235 a_2363_n2734# a_n131_n3054# a_2273_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X236 a_5456_412# a_5402_174# a_5360_46# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X237 a_5360_46# a_3177_n4294# a_5288_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X238 a_6153_n828# B14 a_5402_n1066# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X239 a_541_n2434# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X240 a_1479_n1494# B3 a_1201_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X241 a_1479_n3974# B7 a_1201_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X242 a_3434_n1546# a_3946_n1066# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X243 a_3861_n3080# B8 a_6023_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X244 a_4363_n2068# A9 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X245 a_1467_n3308# A7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X246 DGND B9 a_4000_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 a_3874_n3700# a_5402_n3546# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X248 DVDD B13 a_4000_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 DGND B12 a_5456_46# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X250 a_2569_n4255# a_1968_n4294# a_2497_n4255# DVDD sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X251 a_n41_n4294# a_n71_n4320# a_n131_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X252 a_n41_n4294# B6 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X253 DGND B8 a_5819_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X254 a_n71_n4320# B6 a_315_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X255 a_2569_n1448# a_2315_n1775# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X256 a_2569_n3928# a_2315_n4255# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X257 DVDD B11 a_4363_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X258 a_4697_n3308# B11 a_3946_n3546# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X259 a_1261_n3080# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 DVDD A11 a_4523_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X261 a_n131_n3054# a_n71_n3080# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X262 a_894_n2068# a_143_n2276# a_798_n2434# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X263 a_1291_n1814# B3 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X264 a_1641_46# a_636_n574# a_1557_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X265 DVDD A8 a_5456_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X266 a_2422_n828# B3 a_2350_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X267 DGND a_n131_n1814# a_2543_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X268 a_6023_n3974# A10 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X269 a_6023_n1494# A14 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X270 a_4691_n254# A13 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 a_1641_n828# a_636_n1814# a_1557_n1194# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X272 a_11_n2068# A4 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X273 DVDD A14 a_6153_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X274 DVDD B9 a_4691_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X275 a_2350_n2434# a_636_n3054# a_2254_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X276 a_541_n1194# B2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X277 a_541_n3674# B6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X278 a_6023_n1814# A14 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X279 DVDD A12 a_6153_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X280 a_5360_n1194# a_4204_n574# a_5288_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X281 a_2254_n1194# a_1557_n1194# a_1997_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X282 a_2254_n3674# a_1557_n3674# a_1997_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X283 a_966_n2068# B4 a_894_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X284 DVDD B14 a_5456_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X285 a_5288_n1194# B14 a_5192_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X286 a_5288_n3674# B10 a_5192_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X287 a_3711_n2734# a_3669_n2822# a_3627_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 a_5192_n2068# A8 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X289 a_798_46# a_101_46# a_541_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X290 a_3861_n600# a_5773_n574# a_6023_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X291 a_3832_412# B13 a_3736_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X292 a_6023_n574# A12 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X293 a_4000_412# a_3874_20# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X294 DVDD A5 a_1641_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X295 a_3736_412# A13 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X296 a_2783_n1775# Cin a_2569_n1775# DVDD sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X297 DGND B7 a_1261_n4320# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X298 DGND B3 a_1261_n1840# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X299 DGND A13 a_4000_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X300 a_3543_n2822# a_5773_n4294# a_6023_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X301 a_966_46# B0 a_894_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X302 a_5360_n3674# a_4204_n3054# a_5288_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X303 a_5456_n2434# a_5402_n2306# a_5360_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X304 DVDD a_2273_n254# a_2783_n1775# DVDD sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X305 a_1641_n3308# a_636_n4294# a_1557_n3674# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X306 a_6153_412# B12 a_5402_174# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 a_5773_n3054# B8 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X308 DGND A5 a_2422_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X309 a_2422_n3308# B7 a_2350_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X310 a_541_n1194# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X311 a_541_n3674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X312 a_1291_n1814# a_1261_n1840# a_1201_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X313 a_966_412# B0 a_894_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X314 DGND B13 a_4000_46# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_4441_n574# B13 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_1261_n1840# B3 a_1647_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X317 a_3543_n2822# B10 a_6023_n3974# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X318 a_3543_n342# B14 a_6023_n1494# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X319 a_n71_n600# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 DGND a_101_n2434# a_636_n3054# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X321 DGND B15 a_4000_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X322 DGND B11 a_4000_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X323 a_1467_n2068# A5 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X324 DVDD a_1201_n574# a_2273_n254# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X325 a_2569_n1775# Cin a_2569_n1448# DGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X326 a_2569_n4255# a_143_n2276# a_2569_n3928# DGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X327 a_3627_n2734# a_3543_n2822# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X328 a_185_n2434# a_143_n2276# a_101_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_3322_n1582# a_3765_n600# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X330 DGND a_1557_46# a_143_n1036# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X331 a_1261_n600# B1 a_1647_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X332 DGND B14 a_5819_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X333 DGND B10 a_5819_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X334 a_5402_174# a_3177_n4294# a_5819_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_2783_n4255# a_143_n2276# a_2569_n4255# DVDD sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X336 DVDD B9 a_4363_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X337 a_5192_n828# A14 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X338 a_1261_n4320# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X339 DVDD A5 a_1291_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 a_n131_n1814# a_n71_n1840# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X341 a_1261_n1840# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X342 a_n131_n4294# a_n71_n4320# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X343 a_4697_n2068# B9 a_3946_n2306# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X344 DVDD B14 a_6023_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X345 a_5192_412# A12 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X346 DGND a_n131_n4294# a_2543_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X347 DVDD a_2273_n2734# a_2783_n4255# DVDD sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X348 DVDD a_143_n3516# a_541_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X349 a_1557_n3674# B7 a_1467_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X350 DGND a_2273_n2734# a_2790_n3928# DGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X351 DGND a_2273_n254# a_2790_n1448# DGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X352 a_1641_n3308# B7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X353 a_4000_n3308# a_3874_n3700# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 a_3904_n2434# a_3874_n2460# a_3832_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X355 a_4204_n3054# a_3946_n2306# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X356 a_2350_n3674# a_636_n4294# a_2254_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X357 a_1647_n1814# A3 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X358 a_2350_n1194# a_636_n1814# a_2254_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X359 DVDD B11 a_4691_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X360 a_5288_412# B12 a_5192_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X361 DVDD A11 a_4697_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X362 a_n41_n574# a_n71_n600# a_n131_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X363 a_3226_n1582# a_3177_n4294# a_3368_n1775# DVDD sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X364 a_1997_412# A1 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X365 DVDD A0 a_966_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X366 a_4204_n574# a_3946_174# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X367 DVDD A13 a_4000_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X368 a_1291_n3054# B5 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X369 DVDD A1 a_1291_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X370 a_3322_n1582# a_3543_n342# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X371 a_n41_n574# B0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X372 DVDD a_636_n1814# a_1997_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X373 a_5819_n2434# A8 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X374 DVDD A11 a_4000_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X375 a_5456_n1194# a_5402_n1066# a_5360_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X376 a_5456_n3674# a_5402_n3546# a_5360_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X377 a_5360_n2434# a_2995_n4294# a_5288_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X378 a_1997_46# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X379 a_5402_174# a_3177_n4294# a_5819_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X380 a_1641_n2068# a_636_n3054# a_1557_n2434# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X381 a_5773_n4294# B10 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X382 a_5773_n1814# B14 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X383 DGND Cin a_541_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X384 a_5456_46# a_3177_n4294# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X385 DGND A3 a_2422_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X386 DGND A7 a_2422_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X387 a_2422_n2068# B5 a_2350_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X388 a_2995_n4294# a_2569_n4255# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X389 a_3226_n4062# a_2995_n4294# a_3368_n4255# DVDD sky130_fd_pr__pfet_01v8 ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X390 a_6023_n3054# A8 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X391 DVDD B15 a_4363_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X392 a_143_n2276# a_2569_n1775# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X393 DVDD A12 a_5855_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X394 DGND A1 a_2422_46# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X395 DGND a_101_n1194# a_636_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X396 DGND a_101_n3674# a_636_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X397 a_6153_n2434# B8 a_5402_n2306# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X398 a_1557_46# B1 a_1467_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X399 a_185_n3674# a_143_n3516# a_101_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X400 a_185_n1194# a_143_n1036# a_101_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X401 a_101_46# B0 a_11_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X402 a_5855_n1814# B14 a_5773_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X403 DVDD a_636_n574# a_1997_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X404 a_143_n2276# a_2569_n1775# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X405 a_1201_n574# a_1261_n600# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X406 DVDD A7 a_1291_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 a_4000_n2434# a_3946_n2306# a_3904_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X408 DVDD a_101_n1194# a_636_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X409 a_3795_n2734# a_3765_n3080# a_3711_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X410 DVDD a_143_n2276# a_541_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X411 a_1261_n600# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 a_185_n2434# B4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X413 a_1557_n2434# B5 a_1467_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X414 a_1641_n2068# B5 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X415 a_2908_n600# a_3874_n1220# a_3832_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X416 a_3904_n3674# a_3874_n3700# a_3832_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X417 a_1997_n828# B3 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X418 a_1291_n3054# a_1261_n3080# a_1201_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X419 a_4000_n2068# a_3874_n2460# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X420 a_3434_n4026# a_3946_n3546# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X421 a_1261_n3080# B5 a_1647_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X422 a_2543_n2734# a_1201_n4294# a_2459_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X423 a_894_412# Cin a_798_46# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X424 a_541_n3308# B6 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X425 DGND a_636_n3054# a_1997_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X426 a_101_n2434# B4 a_11_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X427 DVDD A9 a_4697_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.063 ps=0.72 w=0.42 l=0.15
X428 DVDD a_n131_n1814# a_2273_n254# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X429 a_5402_n2306# a_2995_n4294# a_5819_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X430 a_2273_n2734# a_n131_n3054# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X431 a_798_46# a_101_46# a_541_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X432 a_2254_n3674# a_1557_n3674# a_1997_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X433 DGND A8 a_5773_n3054# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X434 a_4691_n574# A13 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X435 DVDD B13 a_4363_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X436 DGND A1 a_1641_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 a_5288_n3308# B10 a_5192_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X438 a_1291_n4294# B7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X439 DVDD B8 a_6023_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X440 a_1641_412# B1 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X441 a_5288_46# B12 a_5192_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X442 DVDD B12 a_5456_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X443 DVDD a_143_n1036# a_541_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X444 DGND A4 a_185_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X445 a_5819_n3674# A10 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 a_5819_n1194# A14 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X447 DVDD A9 a_4000_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X448 a_2363_n254# a_n131_n574# a_2273_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X449 a_1647_n3054# A5 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X450 a_5456_46# a_5402_174# a_5360_46# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X451 a_2459_n2734# a_1201_n3054# a_2363_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X452 a_6023_n4294# A10 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 a_541_n3308# A6 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X454 a_1479_n254# B1 a_1201_n574# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X455 DGND B8 a_5456_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X456 a_3736_n2434# A9 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X457 DVDD B11 a_4000_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X458 a_6153_n1194# B14 a_5402_n1066# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X459 a_6153_n3674# B10 a_5402_n3546# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 DGND A13 a_4697_46# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X461 a_3765_n600# B13 a_4691_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X462 DVDD B10 a_5819_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X463 a_3322_n4062# a_3861_n3080# a_3795_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X464 DGND a_101_46# a_636_n574# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X465 a_4523_n574# B13 a_4441_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X466 a_n71_n3080# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X467 a_315_n574# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X468 DGND B12 a_5819_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X469 a_4000_n1194# a_3946_n1066# a_2908_n600# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X470 a_4000_n3674# a_3946_n3546# a_3904_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X471 DVDD a_3669_n2822# a_3322_n4062# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X472 a_4441_n3054# B9 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X473 DVDD A1 a_1641_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X474 a_1467_n828# A3 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X475 a_185_n1194# B2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X476 a_185_n3674# B6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X477 DVDD B14 a_5819_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X478 DVDD a_1557_46# a_143_n1036# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X479 DGND a_1557_n2434# a_143_n3516# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X480 DGND A8 a_6153_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X481 a_5402_n1066# a_4204_n574# a_5819_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X482 a_1291_n4294# a_1261_n4320# a_1201_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X483 a_3946_n1066# a_3874_n1220# a_4363_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X484 a_1261_n4320# B7 a_1647_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X485 a_2350_n3308# a_636_n4294# a_2254_n3674# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X486 a_5456_n2434# a_2995_n4294# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 a_541_n2068# B4 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X488 DGND a_636_n1814# a_1997_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X489 DGND a_636_n4294# a_1997_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X490 a_101_n3674# B6 a_11_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X491 a_185_n828# B2 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X492 a_3832_n828# B15 a_3736_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X493 a_101_n1194# B2 a_11_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X494 a_5402_n1066# a_4204_n574# a_5819_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X495 a_5402_n3546# a_4204_n3054# a_5819_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 a_3368_n1775# a_3322_n1582# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X497 a_5855_n3054# B8 a_5773_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X498 a_2254_n2434# a_1557_n2434# a_1997_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X499 DGND A10 a_5773_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X500 DGND A14 a_5773_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X501 a_5288_n2068# B8 a_5192_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X502 a_5456_412# a_3177_n4294# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X503 DVDD B10 a_6023_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X504 DVDD a_101_n2434# a_636_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X505 a_3322_n4062# a_3543_n2822# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X506 a_798_n2434# a_101_n2434# a_541_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X507 DGND A2 a_185_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X508 DGND A6 a_185_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 a_2543_n254# a_1201_n1814# a_2459_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 DGND A13 a_4441_n574# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X511 a_1557_n1194# B3 a_1467_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X512 DVDD A14 a_5855_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X513 DGND B0 a_n71_n600# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X514 a_4204_n574# a_3946_174# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X515 a_5456_n3308# a_5402_n3546# a_5360_n3674# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X516 a_1647_n4294# A7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 DGND a_4441_n574# a_3765_n600# DGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X518 a_3832_n2434# B9 a_3736_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X519 a_1997_n2434# B5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X520 DVDD a_n131_n4294# a_2273_n2734# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X521 DVDD A7 a_2422_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X522 a_3368_n4255# a_3322_n4062# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X523 a_3946_n2306# a_3874_n2460# a_4363_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X524 a_541_n2068# A4 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 a_541_46# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X526 DGND B14 a_5456_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X527 a_3736_n3674# A11 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X528 DGND B10 a_5456_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X529 a_3736_n1194# A15 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X530 a_3368_n3928# a_3322_n4062# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X531 a_3368_n1448# a_3322_n1582# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X532 a_5456_n828# a_4204_n574# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X533 DVDD B9 a_4000_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X534 DGND A12 a_6153_46# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X535 a_3861_n600# B12 a_6023_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X536 a_185_n3308# a_143_n3516# a_101_n3674# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X537 DVDD B8 a_5819_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X538 a_185_n828# a_143_n1036# a_101_n1194# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 a_1997_n2434# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X540 DGND B13 a_4363_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X541 DGND a_2908_n600# S15 DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X542 a_n71_n1840# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X543 a_n71_n4320# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X544 DGND A4 a_966_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X545 a_2422_412# B1 a_2350_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X546 a_3589_n3928# a_2995_n4294# a_3226_n4062# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X547 a_4441_n4294# B11 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X548 a_4441_n1814# B15 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X549 a_3589_n1448# a_3177_n4294# a_3226_n1582# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X550 DGND A14 a_6153_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X551 DGND a_1557_n1194# a_1968_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X552 DGND A10 a_6153_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.063 ps=0.72 w=0.42 l=0.15
X553 DGND a_1557_n3674# a_1968_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X554 a_3904_n3674# a_3874_n3700# a_3832_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X555 a_4363_n2434# A9 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X556 DGND A4 a_147_n2734# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X557 a_541_412# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X558 a_5456_n1194# a_4204_n574# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X559 a_5456_n3674# a_4204_n3054# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X560 a_2350_n2068# a_636_n3054# a_2254_n2434# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X561 a_315_n1814# A2 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X562 a_3711_n254# a_3669_n342# a_3627_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X563 a_185_46# Cin a_101_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X564 DGND A0 a_147_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X565 a_4691_n2734# A9 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X566 a_4523_n1814# B15 a_4441_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X567 DVDD A1 a_2422_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X568 a_1647_n574# A1 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X569 a_3669_n342# a_4441_n1814# a_4691_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X570 a_5855_n4294# B10 a_5773_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X571 a_1997_n828# A3 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X572 DVDD a_1557_n1194# a_1968_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X573 a_5819_412# A12 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X574 a_2995_n4294# a_2569_n4255# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X575 DGND A8 a_5456_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06195 ps=0.715 w=0.42 l=0.15
X576 a_894_n2434# a_143_n2276# a_798_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X577 a_1291_n574# a_1261_n600# a_1201_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X578 DVDD A3 a_2422_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X579 a_1641_46# B1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X580 DVDD a_101_n3674# a_636_n4294# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X581 a_3685_n1775# a_3434_n1546# a_3226_n1582# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X582 a_185_46# B0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X583 a_3946_174# a_3874_20# a_4363_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X584 a_798_n1194# a_101_n1194# a_541_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X585 a_798_n3674# a_101_n3674# a_541_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X586 DVDD a_2273_n254# a_2315_n1775# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X587 a_3874_n2460# a_5402_n2306# DGND DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X588 a_11_n2434# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X589 a_5819_n3308# A10 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X590 a_11_412# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1575 ps=1.59 w=0.42 l=0.15
X591 a_101_46# B0 a_11_46# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X592 a_4000_n828# a_3874_n1220# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X593 a_147_n2734# B4 a_n131_n3054# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X594 a_5456_n2068# a_5402_n2306# a_5360_n2434# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X595 a_1997_n1194# B3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X596 a_3832_n1194# B15 a_3736_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X597 a_3832_n3674# B11 a_3736_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X598 a_1997_n3674# B7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X599 DGND B4 a_n71_n3080# DGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X600 a_3226_n4062# a_3434_n4026# a_3368_n3928# DGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X601 a_3226_n1582# a_3434_n1546# a_3368_n1448# DGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X602 a_5456_n828# a_5402_n1066# a_5360_n1194# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X603 DVDD A5 a_2422_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X604 a_3946_n1066# a_3874_n1220# a_4363_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X605 a_3946_n3546# a_3874_n3700# a_4363_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X606 a_3322_n4062# a_3765_n3080# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X607 a_966_n2434# B4 a_894_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X608 DGND A9 a_4441_n3054# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X609 a_4000_n828# a_3946_n1066# a_2908_n600# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X610 a_5192_n2434# A8 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X611 DVDD a_3655_n1516# a_3685_n1775# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X612 DVDD Cin a_541_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X613 a_2273_n254# a_n131_n574# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X614 a_6153_n3308# B10 a_5402_n3546# DVDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
X615 DGND A5 a_1641_n2434# DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X616 a_2273_n2734# a_1201_n4294# DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X617 a_3685_n4255# a_3434_n4026# a_3226_n4062# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X618 a_185_n2068# a_143_n2276# a_101_n2434# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X619 a_1997_n1194# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 a_1997_n3674# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X621 DVDD a_2273_n2734# a_2315_n4255# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X622 a_1291_n574# B1 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X623 DGND a_3655_n3996# a_3589_n3928# DGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X624 DGND a_3655_n1516# a_3589_n1448# DGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X625 a_1997_412# B1 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X626 DVDD B12 a_5819_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X627 DGND a_3226_n4062# a_3177_n4294# DGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X628 DVDD A8 a_5855_n3054# DVDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 DGND a_3226_n1582# a_3177_n1814# DGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X630 DGND a_2273_n254# a_2315_n1775# DGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X631 DGND a_2273_n2734# a_2315_n4255# DGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X632 DVDD A3 a_1641_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X633 DGND A2 a_966_n1194# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X634 DGND A6 a_966_n3674# DGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X635 a_4000_n3308# a_3946_n3546# a_3904_n3674# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X636 a_4000_412# a_3946_174# a_3904_46# DVDD sky130_fd_pr__pfet_01v8 ad=0.06195 pd=0.715 as=0.0693 ps=0.75 w=0.42 l=0.15
X637 a_185_412# B0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X638 a_5819_46# A12 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X639 a_185_n3308# B6 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X640 a_5773_n574# B12 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X641 a_2350_n828# a_636_n1814# a_2254_n1194# DVDD sky130_fd_pr__pfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X642 a_3736_n828# A15 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1575 ps=1.59 w=0.42 l=0.15
X643 DVDD B13 a_4691_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X644 a_4363_n1194# A15 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X645 a_4363_n3674# A11 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X646 a_3904_n2434# a_3874_n2460# a_3832_n2068# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X647 a_3904_46# a_3874_20# a_3832_412# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X648 a_3322_n1582# a_3861_n600# a_3795_n254# DGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X649 DGND A2 a_147_n1494# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X650 DGND A6 a_147_n3974# DGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X651 a_1467_n2434# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.1596 ps=1.6 w=0.42 l=0.15
X652 DVDD A2 a_966_n828# DVDD sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.59 as=0.0693 ps=0.75 w=0.42 l=0.15
X653 DVDD a_101_46# a_636_n574# DVDD sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X654 DVDD a_3655_n3996# a_3685_n4255# DVDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X655 DVDD a_3226_n1582# a_3177_n1814# DVDD sky130_fd_pr__pfet_01v8 ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X656 DVDD a_636_n4294# a_1997_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X657 a_101_n3674# B6 a_11_n3308# DVDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
.ends

