** sch_path: /home/global/EE23B038/tutorial_6/6_1a/tutorial_6_1.sch
**.subckt tutorial_6_1
Vin1 Vin GND PULSE(0 1.8 10ps 5ps 5ps 100ps 250ps)
Vdd1 VDD GND 1.8
x1 VDD Vin Vout GND inv
x2 VDD Vout net1 GND inv
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.include inv_extracted.spice
.control
tran 0.01p 250p
plot v(Vout) v(Vin)
meas tran thl trig v(Vin) val=0.9 rise=1 targ v(Vout) val=0.9 fall=1
meas tran tlh trig v(Vin) val=0.9 fall=1 targ v(Vout) val=0.9 rise=1
let delay = ( $&thl + $&tlh ) / 2
echo delay : $&delay
.endc

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
