* NGSPICE file created from inv.ext - technology: sky130A

.subckt inv in out DVDD DGND
X0 out in DGND DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 out in DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
.ends

