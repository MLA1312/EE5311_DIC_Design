** sch_path: /home/global/EE23B038/tutorial_8/fa16.sch
.subckt fa16 S15 DVDD A12 A13 A14 A15 A9 A8 A10 A11 B13 B12 A6 B14 A5 A4 B15 A7 A2 B11 B10 A0 B9 B8 A1 A3 B6 B5 B4 B7 B2 B0 B3 B1
+ Cin DGND
*.PININFO A0:I B0:I Cin:I A1:I B1:I A2:I B2:I A3:I B3:I A4:I B4:I A5:I B5:I A6:I B6:I A7:I B7:I A8:I B8:I A9:I B9:I A10:I B10:I
*+ A11:I B11:I A12:I B12:I A13:I B13:I A14:I B14:I A15:I B15:I DGND:B DVDD:B S15:O
x1 DVDD DGND A0 B0 Cin net1 net54 fa
x6 DVDD A0 B0 net11 DGND xor2
x2 net1 net3 DVDD DGND inv
x3 DVDD DGND A1 B1 net3 net2 net55 fa
x4 DVDD A1 B1 net10 DGND xor2
x5 net2 net5 DVDD DGND inv
x7 DVDD DGND A2 B2 net5 net4 net56 fa
x8 DVDD A2 B2 net8 DGND xor2
x9 net4 net7 DVDD DGND inv
x10 DVDD DGND A3 B3 net7 net6 net57 fa
x11 DVDD A3 B3 net9 DGND xor2
x12 net6 net13 DVDD DGND inv
x13 DVDD net11 net10 net9 net8 net12 DGND nand4
x14 DVDD net12 Cin net13 C1 DGND mux2
x15 DVDD DGND A4 B4 C1 net14 net58 fa
x16 DVDD A4 B4 net24 DGND xor2
x17 net14 net16 DVDD DGND inv
x18 DVDD DGND A5 B5 net16 net15 net59 fa
x19 DVDD A5 B5 net23 DGND xor2
x20 net15 net18 DVDD DGND inv
x21 DVDD DGND A6 B6 net18 net17 net60 fa
x22 DVDD A6 B6 net21 DGND xor2
x23 net17 net20 DVDD DGND inv
x24 DVDD DGND A7 B7 net20 net19 net61 fa
x25 DVDD A7 B7 net22 DGND xor2
x26 net19 net26 DVDD DGND inv
x27 DVDD net24 net23 net22 net21 net25 DGND nand4
x28 DVDD net25 C1 net26 C2 DGND mux2
x29 DVDD DGND A8 B8 C2 net27 net62 fa
x30 DVDD A8 B8 net37 DGND xor2
x31 net27 net29 DVDD DGND inv
x32 DVDD DGND A9 B9 net29 net28 net63 fa
x33 DVDD A9 B9 net36 DGND xor2
x34 net28 net31 DVDD DGND inv
x35 DVDD DGND A10 B10 net31 net30 net64 fa
x36 DVDD A10 B10 net34 DGND xor2
x37 net30 net33 DVDD DGND inv
x38 DVDD DGND A11 B11 net33 net32 net65 fa
x39 DVDD A11 B11 net35 DGND xor2
x40 net32 net39 DVDD DGND inv
x41 DVDD net37 net36 net35 net34 net38 DGND nand4
x42 DVDD net38 C2 net39 C3 DGND mux2
x43 DVDD DGND A12 B12 C3 net40 net66 fa
x44 DVDD A12 B12 net50 DGND xor2
x45 net40 net42 DVDD DGND inv
x46 DVDD DGND A13 B13 net42 net41 net67 fa
x47 DVDD A13 B13 net49 DGND xor2
x48 net41 net44 DVDD DGND inv
x49 DVDD DGND A14 B14 net44 net43 net68 fa
x50 DVDD A14 B14 net47 DGND xor2
x51 net43 net46 DVDD DGND inv
x52 DVDD DGND A15 B15 net46 net45 net53 fa
x53 DVDD A15 B15 net48 DGND xor2
x54 net45 net52 DVDD DGND inv
x55 DVDD net50 net49 net48 net47 net51 DGND nand4
x56 DVDD net51 C3 net52 net69 DGND mux2
x57 net53 S15 DVDD DGND inv
.ends

* expanding   symbol:  /home/EE23B038/ee5311/tutorial_8/fa.sym # of pins=7
** sym_path: /home/EE23B038/ee5311/tutorial_8/fa.sym
** sch_path: /home/EE23B038/ee5311/tutorial_8/fa.sch
.subckt fa DVDD DGND A B CIN COUTB SUMB
*.PININFO COUTB:O CIN:I DVDD:B DGND:B SUMB:O B:I A:I
XM3 SUMB CIN net4 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM1 net2 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 net1 B net2 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 SUMB CIN net1 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM5 net4 B net3 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM6 net3 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM7 net5 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 net5 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM9 net5 CIN DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 SUMB COUTB net5 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM11 net6 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM12 net6 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM13 net6 CIN DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM14 SUMB COUTB net6 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM15 COUTB CIN net10 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM16 net7 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM17 COUTB B net7 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM18 COUTB CIN net9 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM19 COUTB B net8 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM20 net8 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM21 net9 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM22 net9 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM23 net10 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM24 net10 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends


* expanding   symbol:  /home/EE23B038/ee5311/tutorial_8/xor2.sym # of pins=5
** sym_path: /home/EE23B038/ee5311/tutorial_8/xor2.sym
** sch_path: /home/EE23B038/ee5311/tutorial_8/xor2.sch
.subckt xor2 DVDD A B Y DGND
*.PININFO DVDD:B DGND:B A:I B:I Y:O
XM2 Y net1 net2 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM1 Y net1 DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM3 net1 B net3 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM4 net3 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM5 net1 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM6 net1 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM7 Y B net4 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM8 net4 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM9 net2 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM10 net2 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
.ends


* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/global/EE23B038/tutorial_8/inv.sym
** sch_path: /home/global/EE23B038/tutorial_8/inv.sch
.subckt inv A Y DVDD DGND
*.PININFO Y:O A:I DVDD:B DGND:B
XM2 Y A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM1 Y A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
.ends


* expanding   symbol:  nand4.sym # of pins=7
** sym_path: /home/global/EE23B038/tutorial_8/nand4.sym
** sch_path: /home/global/EE23B038/tutorial_8/nand4.sch
.subckt nand4 DVDD A B C D Y DGND
*.PININFO Y:O A:I DVDD:B DGND:B B:I C:I D:I
XM2 Y B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM1 Y A net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM3 net1 B net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM4 net2 C net3 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM5 net3 D DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM6 Y A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM7 Y C DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM8 Y D DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
.ends


* expanding   symbol:  mux2.sym # of pins=6
** sym_path: /home/global/EE23B038/tutorial_8/mux2.sym
** sch_path: /home/global/EE23B038/tutorial_8/mux2.sch
.subckt mux2 DVDD S A0 A1 Y DGND
*.PININFO DVDD:B DGND:B A0:I A1:I S:I Y:O
XM2 Y net1 DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM1 Y net1 DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM3 net2 S DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 net1 A0 net2 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM5 Sb S DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.00 nf=1 m=1
XM6 Sb S DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM7 net1 A0 net3 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM8 net3 Sb DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM9 net4 Sb DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 net1 A1 net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM11 net1 A1 net5 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
XM12 net5 S DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 m=1
.ends

.end
