** sch_path: /home/global/EE23B038/tutorial_2/tutorial_2_1a (copy 1).sch
**.subckt tutorial_2_1a (copy 1)
XM1 Vin Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vin Vin GND 1.8
**** begin user architecture code

.control
dc Vin 0 1.8 0.01
plot -i(Vin)
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
