** sch_path: /home/EE23B038/ee5311/tutorial_3/tutorial_3_1d.sch
**.subckt tutorial_3_1d
XM2 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vin1 Vin GND 1.8
Vdd1 VDD GND 1.8
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.control
let vds = 0.8
let index = 1
let N = 2
let vals = vector(N)
while index le N
    alter Vdd1 $&vds
    dc Vin1 0 $&vds 0.01
    let vals[index - 1] = abs(vecmin(dc{$&index}.i(Vdd1)))
    let vds = vds + 1
    let index = index + 1
end
let I0 = vals[0]
let I1 = vals[1]
echo I0max: $&I0 I1max: $&I1
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
