* NGSPICE file created from inv.ext - technology: sky130A
.subckt inv DVDD in out DGND
X0 out.t1 in.t0 DGND.t1 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 out.t0 in.t1 DVDD.t1 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
R0 in.n0 in.t1 260.779
R1 in.n0 in.t0 177.232
R2 in in.n0 154.37
R3 DGND DGND.t0 4634.04
R4 DGND DGND.t1 275.918
R5 out out.t0 416.603
R6 out out.t1 271.904
R7 DVDD DVDD.t0 949.298
R8 DVDD DVDD.t1 398.106
C0 out DVDD 0.103082f
C1 in DVDD 0.104904f
C2 out in 0.039201f
C3 out DGND 0.12215f
C4 in DGND 0.227683f
C5 DVDD DGND 0.773835f
.ends
