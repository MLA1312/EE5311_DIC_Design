* NGSPICE file created from nors.ext - technology: sky130A
.subckt nors DVDD Y A DGND
X0 a_924_288# Y.t8 DGND.t19 DGND.t18 sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.126 ps=1.44 w=0.42 l=0.15
X1 DGND.t1 A.t0 Y.t5 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.105 ps=0.92 w=0.42 l=0.15
X2 Y.t4 DGND.t13 DGND.t15 DGND.t14 sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.126 ps=1.44 w=0.42 l=0.15
X3 DGND.t12 DGND.t10 Y.t6 DGND.t11 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.105 ps=0.92 w=0.42 l=0.15
X4 a_834_288# DGND.t20 DVDD.t19 DVDD.t18 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X5 a_924_288# Y.t9 a_834_288# DVDD.t23 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X6 DGND.t17 Y.t10 a_924_288# DGND.t16 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.105 ps=0.92 w=0.42 l=0.15
X7 DVDD.t17 DGND.t21 a_834_288# DVDD.t16 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X8 Y.t7 A.t1 DGND.t3 DGND.t2 sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.126 ps=1.44 w=0.42 l=0.15
X9 a_834_288# DGND.t22 DVDD.t15 DVDD.t14 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X10 a_834_288# Y.t11 a_924_288# DVDD.t22 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X11 DVDD.t13 DGND.t23 a_n702_288# DVDD.t12 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X12 DVDD.t11 DGND.t24 a_834_288# DVDD.t10 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X13 a_924_288# Y.t12 a_834_288# DVDD.t21 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X14 a_n702_288# DGND.t25 DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X15 a_924_288# DGND.t7 DGND.t9 DGND.t8 sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.126 ps=1.44 w=0.42 l=0.15
X16 Y.t0 A.t2 a_n702_288# DVDD.t3 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X17 a_834_288# Y.t13 a_924_288# DVDD.t20 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X18 DVDD.t7 DGND.t26 a_n702_288# DVDD.t6 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X19 DGND.t6 DGND.t4 a_924_288# DGND.t5 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.105 ps=0.92 w=0.42 l=0.15
X20 a_n702_288# A.t3 Y.t1 DVDD.t2 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X21 a_n702_288# DGND.t27 DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X22 Y.t2 A.t4 a_n702_288# DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X23 a_n702_288# A.t5 Y.t3 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
R0 Y.n10 Y.n9 1019.94
R1 Y.n2 Y.n1 422.231
R2 Y.n5 Y.t9 383.522
R3 Y.n2 Y.n0 324.348
R4 Y.n11 Y.n10 229.648
R5 Y.n11 Y.n3 219.636
R6 Y.n10 Y.n4 215.871
R7 Y.n9 Y.n8 202.13
R8 Y.n7 Y.t11 199.227
R9 Y.n6 Y.t12 199.227
R10 Y.n5 Y.t13 199.227
R11 Y.n7 Y.n6 184.294
R12 Y.n6 Y.n5 184.294
R13 Y Y.n2 177.695
R14 Y Y.n11 173.177
R15 Y.n8 Y.n7 149.421
R16 Y.n8 Y.t10 91.5805
R17 Y.n9 Y.t8 91.5805
R18 Y.n3 Y.t5 71.4291
R19 Y.n3 Y.t7 71.4291
R20 Y.n4 Y.t6 71.4291
R21 Y.n4 Y.t4 71.4291
R22 Y.n0 Y.t3 58.6315
R23 Y.n0 Y.t2 58.6315
R24 Y.n1 Y.t1 58.6315
R25 Y.n1 Y.t0 58.6315
R26 DGND.t11 DGND.t18 11334.6
R27 DGND.n18 DGND.t8 3417.48
R28 DGND.t16 DGND.n18 3417.48
R29 DGND.n19 DGND.t14 3417.48
R30 DGND.n19 DGND.t0 3417.48
R31 DGND.t8 DGND.t5 1851.13
R32 DGND.t18 DGND.t16 1851.13
R33 DGND.t14 DGND.t11 1851.13
R34 DGND.t0 DGND.t2 1851.13
R35 DGND.n20 DGND.n19 1216.38
R36 DGND.n18 DGND.n17 1216.38
R37 DGND.n8 DGND.t27 383.522
R38 DGND.n1 DGND.t20 383.522
R39 DGND.n11 DGND.t10 287.392
R40 DGND.n4 DGND.t4 287.392
R41 DGND DGND.t3 261.031
R42 DGND.n21 DGND.t1 260.805
R43 DGND.n15 DGND.t19 260.805
R44 DGND.n16 DGND.t17 260.805
R45 DGND.n6 DGND.t6 259.818
R46 DGND.n0 DGND.t15 259.675
R47 DGND.n14 DGND.t12 259.675
R48 DGND.n7 DGND.t9 259.675
R49 DGND.n10 DGND.t26 199.227
R50 DGND.n8 DGND.t23 199.227
R51 DGND.n9 DGND.t25 199.227
R52 DGND.n3 DGND.t24 199.227
R53 DGND.n1 DGND.t21 199.227
R54 DGND.n2 DGND.t22 199.227
R55 DGND.n9 DGND.n8 184.294
R56 DGND.n10 DGND.n9 184.294
R57 DGND.n2 DGND.n1 184.294
R58 DGND.n3 DGND.n2 184.294
R59 DGND.n12 DGND.t10 176.198
R60 DGND.n5 DGND.t4 175.305
R61 DGND.n5 DGND.t7 175.305
R62 DGND.n12 DGND.t13 174.413
R63 DGND.n13 DGND.n12 161.3
R64 DGND.n6 DGND.n5 161.3
R65 DGND.n11 DGND.n10 131.748
R66 DGND.n4 DGND.n3 131.748
R67 DGND.t13 DGND.n11 91.5805
R68 DGND.t7 DGND.n4 91.5805
R69 DGND.n15 DGND.n14 0.919771
R70 DGND.n16 DGND.n15 0.286958
R71 DGND.n17 DGND.n7 0.254406
R72 DGND.n17 DGND.n16 0.254406
R73 DGND.n20 DGND.n0 0.254406
R74 DGND.n21 DGND.n20 0.254406
R75 DGND.n14 DGND.n13 0.145031
R76 DGND.n7 DGND.n6 0.143729
R77 DGND.n13 DGND.n0 0.142427
R78 DGND DGND.n21 0.0603958
R79 A A.t3 527.254
R80 A.n1 A.t4 383.522
R81 A.n0 A.t1 293.709
R82 A.n2 A.t2 199.227
R83 A.n1 A.t5 199.227
R84 A.t3 A.n3 199.227
R85 A.n3 A.n2 184.294
R86 A.n2 A.n1 184.294
R87 A.n3 A.n0 149.421
R88 A.n0 A.t0 91.5805
R89 DVDD.t4 DVDD.t23 809.26
R90 DVDD.n8 DVDD.t10 703.705
R91 DVDD.t22 DVDD.n8 703.705
R92 DVDD.n9 DVDD.t6 703.705
R93 DVDD.n9 DVDD.t2 703.705
R94 DVDD.t16 DVDD.t18 381.173
R95 DVDD.t14 DVDD.t16 381.173
R96 DVDD.t10 DVDD.t14 381.173
R97 DVDD.t21 DVDD.t22 381.173
R98 DVDD.t20 DVDD.t21 381.173
R99 DVDD.t23 DVDD.t20 381.173
R100 DVDD.t12 DVDD.t4 381.173
R101 DVDD.t8 DVDD.t12 381.173
R102 DVDD.t6 DVDD.t8 381.173
R103 DVDD.t2 DVDD.t3 381.173
R104 DVDD.t3 DVDD.t0 381.173
R105 DVDD.t0 DVDD.t1 381.173
R106 DVDD.n2 DVDD.n1 372.507
R107 DVDD.n2 DVDD.n0 372.507
R108 DVDD.n6 DVDD.n5 372.507
R109 DVDD.n6 DVDD.n4 372.507
R110 DVDD DVDD.n9 239.132
R111 DVDD.n8 DVDD.n7 238.904
R112 DVDD.n1 DVDD.t9 58.6315
R113 DVDD.n1 DVDD.t7 58.6315
R114 DVDD.n0 DVDD.t5 58.6315
R115 DVDD.n0 DVDD.t13 58.6315
R116 DVDD.n5 DVDD.t15 58.6315
R117 DVDD.n5 DVDD.t11 58.6315
R118 DVDD.n4 DVDD.t19 58.6315
R119 DVDD.n4 DVDD.t17 58.6315
R120 DVDD.n7 DVDD.n6 9.86691
R121 DVDD.n3 DVDD.n2 9.3005
R122 DVDD.n7 DVDD.n3 1.43409
R123 DVDD DVDD.n3 0.33774
C0 a_834_288# DVDD 0.511125f
C1 Y DVDD 0.540706f
C2 DVDD a_n702_288# 0.50928f
C3 A DVDD 0.422505f
C4 Y a_834_288# 0.103268f
C5 Y a_n702_288# 0.733234f
C6 DVDD a_924_288# 0.238604f
C7 Y A 0.125446f
C8 A a_n702_288# 0.112096f
C9 a_834_288# a_924_288# 0.639339f
C10 Y a_924_288# 0.169494f
C11 a_924_288# a_n702_288# 0.05021f
C12 A a_924_288# 6.13e-20
C13 Y DGND 1.59213f
C14 A DGND 0.557556f
C15 DVDD DGND 4.69206f
C16 a_924_288# DGND 0.631005f
C17 a_834_288# DGND 0.365978f
C18 a_n702_288# DGND 0.258131f
.ends
