** sch_path: /home/EE23B038/ee5311/tutorial_1/nfetsat.sch
**.subckt nfetsat
XM1 net1 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W='0.42 * 1 ' nf=1 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=1
+ m=1
V1 net1 GND 1.8
**** begin user architecture code

.control
set filetype=ascii
dc V1 0 1.8 0.01
wrdata nMOS_ids_vgs.txt -I(V1)
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
